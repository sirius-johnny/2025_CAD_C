VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

USEMINSPACING OBS OFF ;


PROPERTYDEFINITIONS 
LAYER LEF58_CUTCLASS STRING ;
LAYER LEF58_TYPE STRING ;
LAYER LEF58_ENCLOSURE STRING ;
LAYER LEF58_SPACING STRING ;
LAYER LEF58_SPACINGTABLE STRING ;
LAYER LEF58_WIDTH STRING ;
LAYER LEF58_EOLKEEPOUT STRING ;
LAYER LEF58_WIDTHTABLE STRING ; 
LAYER LEF58_RIGHTWAYONGRIDONLY STRING ; 
LAYER LEF58_CORNERSPACING STRING ;
LAYER LEF58_PITCH STRING ;
LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS
LAYER nwell

	TYPE MASTERSLICE ;
	PROPERTY LEF58_TYPE "TYPE NWELL ; " ;
END nwell

LAYER pwell

	TYPE MASTERSLICE ;
	PROPERTY LEF58_TYPE "TYPE PWELL ; " ;
END pwell

LAYER Gate

	TYPE MASTERSLICE ;
END Gate

LAYER Active

	TYPE MASTERSLICE ;
END Active

LAYER V0

	TYPE CUT ;
	SPACING 0.018  ;
	
	WIDTH 0.018 ;
END V0

LAYER M1

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.036 ;
	WIDTH 0.018 ;
	OFFSET 0.0 ;
	AREA 0.000666 ;
	
	SPACING 0.018  ;
	SPACING 0.018 
		RANGE 0.036 1.0  ;
	
	WIREEXTENSION 0.009 ;
	MINWIDTH 0.018 ;
	PROPERTY LEF58_EOLKEEPOUT
	"EOLKEEPOUT 0.018 EXTENSION 0.0 0.0 0.031 ;
	 " ;
	PROPERTY LEF58_CORNERSPACING
	"CORNERSPACING CONVEXCORNER CORNERONLY 0.01 
	WIDTH 0.018 SPACING 0.018 ;
	 " ;
END M1

LAYER V1

	TYPE CUT ;
	SPACING 0.018  ;
	
	WIDTH 0.018 ;
END V1

LAYER M2

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PROPERTY LEF58_PITCH 
	"PITCH  0.036 FIRSTLASTPITCH 0.045 ;" ;
	PITCH 0.036 ;
	WIDTH 0.018 ;
	OFFSET -0.27 ;
	PROPERTY LEF58_RECTONLY 
	"RECTONLY ;" ;
	PROPERTY LEF58_WIDTHTABLE
	"WIDTHTABLE 
    0.018 0.09 0.162 
    0.234 0.306 0.378 ;" ;

	AREA 0.000666 ;
	
	MINSIZE  0.018 0.037  ;
	
	SPACING 0.018  ;
	
	PROPERTY LEF58_SPACING
	"SPACING 0.018 
		ENDOFLINE 0.025 WITHIN 0.02 
			ENDTOEND 0.031 
			PARALLELEDGE 0.025 WITHIN 0.02 ;
	 " ;
	WIREEXTENSION 0.009 ;
	MINWIDTH 0.018 ;
	PROPERTY LEF58_EOLKEEPOUT
	"EOLKEEPOUT 0.025 EXTENSION 0.0 0.013 0.031 CORNERONLY ;
	 " ;
	PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
	PROPERTY LEF58_CORNERSPACING
	"CORNERSPACING CONVEXCORNER
	WIDTH 0.0 SPACING 0.02 ;
	 " ;
END M2

LAYER V2

	TYPE CUT ;
	SPACING 0.018  ;
	
	WIDTH 0.018 ;
END V2

LAYER M3

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.036 ;
	WIDTH 0.018 ;
	OFFSET 0.0 ;
	PROPERTY LEF58_RECTONLY 
	"RECTONLY ;" ;
	PROPERTY LEF58_WIDTHTABLE
	"WIDTHTABLE 
    0.018 0.09 0.162 
    0.234 0.306 0.378 ;" ;

	AREA 0.000666 ;
	
	MINSIZE  0.018 0.037  ;
	
	SPACING 0.018  ;
	
	PROPERTY LEF58_SPACING
	"SPACING 0.018 
		ENDOFLINE 0.025 WITHIN 0.013 
			ENDTOEND 0.031 
			PARALLELEDGE 0.025 WITHIN 0.02 ;
	 " ;
	WIREEXTENSION 0.009 ;
	MINWIDTH 0.018 ;
	PROPERTY LEF58_EOLKEEPOUT
	"EOLKEEPOUT 0.025 EXTENSION 0.0 0.013 0.031 CORNERONLY ;
	 " ;
	PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
	PROPERTY LEF58_CORNERSPACING
	"CORNERSPACING CONVEXCORNER
	WIDTH 0.0 SPACING 0.02 ;
	 " ;
END M3

LAYER V3

	TYPE CUT ;
	PROPERTY LEF58_CUTCLASS
	"CUTCLASS V3_0p864 WIDTH 0.018 LENGTH 0.216 CUTS 8 ;
	CUTCLASS V3_0p480 WIDTH 0.018 LENGTH 0.12 CUTS 4 ;
	CUTCLASS V3 WIDTH 0.018 LENGTH 0.024 ;
	" ;
	PROPERTY LEF58_SPACINGTABLE 
	"SPACINGTABLE		CUTCLASS	      V3	 	V3_0p480	 	V3_0p864	 
	      V3	 	0.034 0.034	0.034 0.034	0.034 0.034
	V3_0p480	 	0.034 0.034	0.034 0.034	0.034 0.034
	V3_0p864	 	0.034 0.034	0.034 0.034	0.034 0.034
 ;
 " ;
	PROPERTY LEF58_ENCLOSURE
	"ENCLOSURE  CUTCLASS V3_0p864  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS V3_0p480  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS V3  ABOVE  EOL 0.024 0.011 0.0 ;
	ENCLOSURE  CUTCLASS V3  BELOW  0.0 0.005  ;
	 " ;
END V3

LAYER M4

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.048 ;
	WIDTH 0.024 ;
	OFFSET 0.003 ;
	PROPERTY LEF58_RECTONLY 
	"RECTONLY ;" ;
	PROPERTY LEF58_WIDTHTABLE
	"WIDTHTABLE 
    0.024 0.12 0.216 
    0.312 0.408 ;" ;

	AREA 0.002 ;
	
	SPACING 0.024  ;
	
	PROPERTY LEF58_SPACING
	"SPACING 0.024 
		ENDOFLINE 0.025 WITHIN 0.04 
			ENDTOEND 0.04  ;
	 " ;
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.024 
		WIDTH 0.025	           		  0.072 ;

	WIREEXTENSION 0.012 ;
	MINWIDTH 0.024 ;
	PROPERTY LEF58_EOLKEEPOUT
	"EOLKEEPOUT 0.025 EXTENSION 0.048 0.024 0.048 CORNERONLY ;
	 " ;
	PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
	PROPERTY LEF58_CORNERSPACING
	"CORNERSPACING CONVEXCORNER CORNERONLY 0.048 
	WIDTH 0.0 SPACING 0.04 ;
	 " ;
END M4

LAYER V4

	TYPE CUT ;
	PROPERTY LEF58_CUTCLASS
	"CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.408 CUTS 16 ;
	CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.312 CUTS 12 ;
	CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.216 CUTS 8 ;
	CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.12 CUTS 4 ;
	CUTCLASS Vx WIDTH 0.024 ;
	" ;
	PROPERTY LEF58_SPACINGTABLE 
	"SPACINGTABLE		CUTCLASS	      Vx	 	Vx_0p480	 	Vx_0p864	 	Vx_1p248	 	Vx_1p632	 
	      Vx	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_0p480	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_0p864	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_1p248	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_1p632	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
 ;
 " ;
	PROPERTY LEF58_ENCLOSURE
	"ENCLOSURE  CUTCLASS Vx_1p632  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_1p248  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_0p864  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_0p480  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx  0.011 0.011  ;
	ENCLOSURE  CUTCLASS Vx  0.0 0.011  ;
	 " ;
END V4

LAYER M5

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.048 ;
	WIDTH 0.024 ;
	OFFSET 0.0 ;
	PROPERTY LEF58_RECTONLY 
	"RECTONLY ;" ;
	PROPERTY LEF58_WIDTHTABLE
	"WIDTHTABLE 
    0.024 0.12 0.216 
    0.312 0.408 0.504 
    0.6 0.696 0.792 
    0.888 0.984 ;" ;

	AREA 0.002 ;
	
	SPACING 0.024  ;
	
	PROPERTY LEF58_SPACING
	"SPACING 0.024 
		ENDOFLINE 0.025 WITHIN 0.04 
			ENDTOEND 0.04  ;
	 " ;
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.024 
		WIDTH 0.025	           		  0.072 ;

	WIREEXTENSION 0.012 ;
	MINWIDTH 0.024 ;
	PROPERTY LEF58_EOLKEEPOUT
	"EOLKEEPOUT 0.025 EXTENSION 0.048 0.024 0.048 CORNERONLY ;
	 " ;
	PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
	PROPERTY LEF58_CORNERSPACING
	"CORNERSPACING CONVEXCORNER CORNERONLY 0.048 
	WIDTH 0.0 SPACING 0.04 ;
	 " ;
	MINIMUMDENSITY 15.0 ;
	MAXIMUMDENSITY 90.0 ;
	DENSITYCHECKWINDOW 20.0 20.0 ;
	DENSITYCHECKSTEP 10.0 ;
END M5

LAYER V5

	TYPE CUT ;
	PROPERTY LEF58_CUTCLASS
	"CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.544 CUTS 16 ;
	CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.416 CUTS 12 ;
	CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.288 CUTS 8 ;
	CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.16 CUTS 4 ;
	CUTCLASS Vx WIDTH 0.024 LENGTH 0.032 ;
	" ;
	PROPERTY LEF58_SPACINGTABLE 
	"SPACINGTABLE		CUTCLASS	      Vx	 	Vx_0p480	 	Vx_0p864	 	Vx_1p248	 	Vx_1p632	 
	      Vx	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_0p480	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_0p864	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_1p248	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_1p632	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
 ;
 " ;
	PROPERTY LEF58_ENCLOSURE
	"ENCLOSURE  CUTCLASS Vx_1p632  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_1p248  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_0p864  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_0p480  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx  EOL 0.024 0.011 0.011 ;
	 " ;
END V5

LAYER M6

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.064 ;
	WIDTH 0.032 ;
	PROPERTY LEF58_RECTONLY 
	"RECTONLY ;" ;
	PROPERTY LEF58_WIDTHTABLE
	"WIDTHTABLE 
    0.032 0.16 0.288 
    0.416 0.544 ;" ;

	AREA 0.0021875 ;
	
	SPACING 0.032  ;
	
	PROPERTY LEF58_SPACING
	"SPACING 0.032 
		ENDOFLINE 0.038 WITHIN 0.04 
			ENDTOEND 0.04  ;
	 " ;
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.032 
		WIDTH 0.033	           		  0.072 ;

	WIREEXTENSION 0.016 ;
	MINWIDTH 0.032 ;
	PROPERTY LEF58_EOLKEEPOUT
	"EOLKEEPOUT 0.05 EXTENSION 0.048 0.032 0.048 CORNERONLY ;
	 " ;
	PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
	PROPERTY LEF58_CORNERSPACING
	"CORNERSPACING CONVEXCORNER CORNERONLY 0.048 
	WIDTH 0.0 SPACING 0.04 ;
	 " ;
END M6

LAYER V6

	TYPE CUT ;
	PROPERTY LEF58_CUTCLASS
	"CUTCLASS Vx_2p176 WIDTH 0.032 LENGTH 0.544 CUTS 16 ;
	CUTCLASS Vx_1p664 WIDTH 0.032 LENGTH 0.416 CUTS 12 ;
	CUTCLASS Vx_1p152 WIDTH 0.032 LENGTH 0.288 CUTS 8 ;
	CUTCLASS Vx_0p640 WIDTH 0.032 LENGTH 0.16 CUTS 4 ;
	CUTCLASS Vx WIDTH 0.032 ;
	" ;
	PROPERTY LEF58_SPACINGTABLE 
	"SPACINGTABLE		CUTCLASS	      Vx	 	Vx_0p640	 	Vx_1p152	 	Vx_1p664	 	Vx_2p176	 
	      Vx	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_0p640	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_1p152	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_1p664	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
	Vx_2p176	 	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034	0.034 0.034
 ;
 " ;
	PROPERTY LEF58_ENCLOSURE
	"ENCLOSURE  CUTCLASS Vx_2p176  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_1p664  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_1p152  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx_0p640  END 0.0 SIDE 0.0  ;
	ENCLOSURE  CUTCLASS Vx  0.011 0.011  ;
	ENCLOSURE  CUTCLASS Vx  0.0 0.011  ;
	 " ;
END V6

LAYER M7

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.064 ;
	WIDTH 0.032 ;
	PROPERTY LEF58_RECTONLY 
	"RECTONLY ;" ;
	PROPERTY LEF58_WIDTHTABLE
	"WIDTHTABLE 
    0.032 0.16 0.288 
    0.416 0.544 ;" ;

	AREA 0.0021875 ;
	
	SPACING 0.032  ;
	
	PROPERTY LEF58_SPACING
	"SPACING 0.03 
		ENDOFLINE 0.038 WITHIN 0.04 
			ENDTOEND 0.04  ;
	 " ;
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.032 
		WIDTH 0.033	           		  0.072 ;

	WIREEXTENSION 0.016 ;
	MINWIDTH 0.032 ;
	PROPERTY LEF58_EOLKEEPOUT
	"EOLKEEPOUT 0.05 EXTENSION 0.048 0.032 0.048 CORNERONLY ;
	 " ;
	PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
	PROPERTY LEF58_CORNERSPACING
	"CORNERSPACING CONVEXCORNER CORNERONLY 0.075 
	WIDTH 0.0 SPACING 0.04 ;
	 " ;
END M7

LAYER V7

	TYPE CUT ;
	SPACING 0.046  ;
	
	WIDTH 0.032 ;
END V7

LAYER M8

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.08 ;
	WIDTH 0.04 ;
	AREA 0.00752 ;
	
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 0.4 1.2 1.8 
		WIDTH 0.0	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.06	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.08	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.12	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.5	           		  0.04 0.04 0.04 0.5 
		WIDTH 1.0	           		  0.04 0.04 0.04 1.0 ;

	WIREEXTENSION 0.02 ;
	MINIMUMCUT 2 WIDTH 1.805 WITHIN 1.705  FROMBELOW  ;
	MINIMUMCUT 2 WIDTH 1.805 WITHIN 1.705  FROMABOVE  ;
	
	MAXWIDTH 2.0 ;
	MINWIDTH 0.04 ;
	MINSTEP 0.04 STEP  ;
	
END M8

LAYER V8

	TYPE CUT ;
	SPACING 0.057  ;
	
	WIDTH 0.04 ;
END V8

LAYER M9

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.08 ;
	WIDTH 0.04 ;
	AREA 0.00752 ;
	
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 0.4 1.2 1.8 
		WIDTH 0.0	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.06	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.08	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.12	           		  0.04 0.04 0.04 0.04 
		WIDTH 0.5	           		  0.04 0.04 0.04 0.5 
		WIDTH 1.0	           		  0.04 0.04 0.04 1.0 ;

	WIREEXTENSION 0.02 ;
	MINIMUMCUT 2 WIDTH 1.805 WITHIN 1.705  FROMABOVE  ;
	
	MINWIDTH 0.04 ;
	MINSTEP 0.04 STEP  ;
	
END M9

LAYER V9

	TYPE CUT ;
	SPACING 0.057  ;
	
	WIDTH 0.04 ;
END V9

LAYER Pad

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.08 ;
	WIDTH 0.04 ;
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 12.0 
		WIDTH 0.0	           		  2.0 2.0 
		WIDTH 12.0	           		  2.0 3.0 ;

	WIREEXTENSION 0.02 ;
	MINIMUMCUT 1 WIDTH 0.04 WITHIN 1.705  FROMBELOW  ;
	MINIMUMCUT 1 WIDTH 0.36 WITHIN 1.705  FROMBELOW  ;
	MINIMUMCUT 2 WIDTH 1.805 WITHIN 1.705  FROMBELOW  ;
	
	MINWIDTH 0.04 ;
	MINIMUMDENSITY 20.0 ;
	MAXIMUMDENSITY 80.0 ;
	DENSITYCHECKWINDOW 100.0 100.0 ;
	DENSITYCHECKSTEP 50.0 ;
END Pad

VIARULE Pad_M9 GENERATE DEFAULT 
	LAYER M9 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER Pad ;
		ENCLOSURE 0.011 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER V9 ;
		RECT -0.016 -0.016 0.016 0.016 ;
		SPACING 0.078 BY 0.078 ;

END Pad_M9 

VIARULE M9_M8 GENERATE DEFAULT 
	LAYER M8 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M9 ;
		ENCLOSURE 0.0 0.02 ;
		WIDTH 0 TO 1000 ;
	LAYER V8 ;
		RECT -0.02 -0.02 0.02 0.02 ;
		SPACING 0.097 BY 0.097 ;

END M9_M8 

VIARULE M8_M7 GENERATE DEFAULT 
	LAYER M7 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M8 ;
		ENCLOSURE 0.011 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER V7 ;
		RECT -0.016 -0.016 0.016 0.016 ;
		SPACING 0.078 BY 0.078 ;

END M8_M7 

VIARULE M7_M6 GENERATE DEFAULT 
	LAYER M6 ;
		ENCLOSURE 0.011 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M7 ;
		ENCLOSURE 0.0 0.011 ;
		WIDTH 0 TO 1000 ;
	LAYER V6 ;
		RECT -0.016 -0.016 0.016 0.016 ;
		SPACING 0.078 BY 0.078 ;

END M7_M6 

VIARULE M6_M5 GENERATE DEFAULT 
	LAYER M5 ;
		ENCLOSURE 0.011 0.0 ;
		WIDTH 0.024 TO 0.024 ;
	LAYER M6 ;
		ENCLOSURE 0.011 0.0 ;
		WIDTH 0.032 TO 0.032 ;
	LAYER V5 ;
		RECT -0.012 -0.016 0.012 0.016 ;
		SPACING 0.058 BY 0.308 ;

END M6_M5 

VIARULE M3_M2widePWR0p936 GENERATE 
	LAYER M2 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M3 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0.234 TO 0.234 ;
	LAYER V2 ;
		RECT -0.117 -0.009 0.117 0.009 ;
		SPACING 0.277 BY 0.036 ;

END M3_M2widePWR0p936 

VIARULE M4_M3widePWR0p864 GENERATE 
	LAYER M3 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0.234 TO 0.234 ;
	LAYER M4 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0.216 TO 0.217 ;
	LAYER V3 ;
		RECT -0.009 -0.108 0.009 0.108 ;
		SPACING 0.036 BY 0.277 ;

END M4_M3widePWR0p864 

VIARULE M5_M4widePWR0p864 GENERATE 
	LAYER M4 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M5 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0.216 TO 0.216 ;
	LAYER V4 ;
		RECT -0.108 -0.012 0.108 0.012 ;
		SPACING 0.532 BY 0.096 ;

END M5_M4widePWR0p864 

VIARULE M6_M5widePWR1p152 GENERATE 
	LAYER M5 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M6 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0.288 TO 0.288 ;
	LAYER V5 ;
		RECT -0.012 -0.144 0.012 0.144 ;
		SPACING 0.096 BY 0.382 ;

END M6_M5widePWR1p152 

VIARULE M7_M6widePWR1p152 GENERATE 
	LAYER M6 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M7 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0.288 TO 0.288 ;
	LAYER V6 ;
		RECT -0.144 -0.016 0.144 0.016 ;
		SPACING 0.532 BY 0.096 ;

END M7_M6widePWR1p152 

VIARULE M2_M1 GENERATE DEFAULT 
	LAYER M1 ;
		ENCLOSURE 0.0 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER M2 ;
		ENCLOSURE 0.002 0.0 ;
		WIDTH 0 TO 1000 ;
	LAYER V1 ;
		RECT -0.009 -0.009 0.009 0.009 ;
		SPACING 0.036 BY 0.036 ;

END M2_M1 

VIA VIA12 DEFAULT 
	LAYER M1 ;
		RECT -0.009 -0.011 0.009 0.011 ;
	LAYER V1 ;
		RECT -0.009 -0.009 0.009 0.009 ;
	LAYER M2 ;
		RECT -0.014 -0.009 0.014 0.009 ;

END VIA12 

VIA VIA23 DEFAULT 
	LAYER M2 ;
		RECT -0.014 -0.009 0.014 0.009 ;
	LAYER V2 ;
		RECT -0.009 -0.009 0.009 0.009 ;
	LAYER M3 ;
		RECT -0.009 -0.014 0.009 0.014 ;

END VIA23 

VIA VIA34 DEFAULT 
	LAYER M3 ;
		RECT -0.009 -0.017 0.009 0.017 ;
	LAYER V3 ;
		RECT -0.009 -0.012 0.009 0.012 ;
	LAYER M4 ;
		RECT -0.02 -0.012 0.02 0.012 ;

END VIA34 

VIA VIA45 DEFAULT 
	LAYER M4 ;
		RECT -0.023 -0.012 0.023 0.012 ;
	LAYER V4 ;
		RECT -0.012 -0.012 0.012 0.012 ;
	LAYER M5 ;
		RECT -0.012 -0.023 0.012 0.023 ;

END VIA45 

VIA VIA56 DEFAULT 
	LAYER M5 ;
		RECT -0.012 -0.027 0.012 0.027 ;
	LAYER V5 ;
		RECT -0.012 -0.016 0.012 0.016 ;
	LAYER M6 ;
		RECT -0.023 -0.016 0.023 0.016 ;

END VIA56 

VIA VIA67 DEFAULT 
	LAYER M6 ;
		RECT -0.027 -0.016 0.027 0.016 ;
	LAYER V6 ;
		RECT -0.016 -0.016 0.016 0.016 ;
	LAYER M7 ;
		RECT -0.016 -0.027 0.016 0.027 ;

END VIA67 

VIA VIA78 DEFAULT 
	LAYER M7 ;
		RECT -0.016 -0.027 0.016 0.027 ;
	LAYER V7 ;
		RECT -0.016 -0.016 0.016 0.016 ;
	LAYER M8 ;
		RECT -0.027 -0.02 0.027 0.02 ;

END VIA78 

VIA VIA89 DEFAULT 
	LAYER M8 ;
		RECT -0.02 -0.02 0.02 0.02 ;
	LAYER V8 ;
		RECT -0.02 -0.02 0.02 0.02 ;
	LAYER M9 ;
		RECT -0.02 -0.02 0.02 0.02 ;

END VIA89 

VIA VIA9Pad DEFAULT 
	LAYER M9 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER V9 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER Pad ;
		RECT -0.05 -0.05 0.05 0.05 ;

END VIA9Pad 

SITE asap7sc7p5t 
	CLASS CORE ;
	SYMMETRY Y ;
	SIZE 0.054 BY 0.27 ;
END asap7sc7p5t 

MACRO A2O1A1Ixp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN A2O1A1Ixp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.214 0.215 0.306 0.233 ;
			RECT 0.288 0.037 0.306 0.233 ;
			RECT 0.262 0.037 0.306 0.055 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.081 0.252 0.19 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.23 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END A2O1A1Ixp33_ASAP7_75t_R

MACRO A2O1A1O1Ixp25_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN A2O1A1O1Ixp25_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.423 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.261 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.127 0.414 0.145 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.207 0.225 0.387 0.243 ;
			RECT 0.04 0.027 0.225 0.045 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END A2O1A1O1Ixp25_ASAP7_75t_R

MACRO AND2x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND2x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.207 0.027 0.306 0.045 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.027 0.18 0.243 ;
			RECT 0.162 0.126 0.203 0.144 ;
			RECT 0.07 0.027 0.088 0.086 ;
			RECT 0.07 0.027 0.18 0.045 ;

	END

END AND2x2_ASAP7_75t_R

MACRO AND2x4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND2x4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.31 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.028 0.252 0.15 ;
			RECT 0.072 0.028 0.252 0.046 ;
			RECT 0.072 0.028 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.107 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.231 0.243 ;
			RECT 0.18 0.064 0.198 0.243 ;
			RECT 0.179 0.182 0.306 0.2 ;
			RECT 0.288 0.121 0.306 0.2 ;
			RECT 0.115 0.064 0.198 0.082 ;

	END

END AND2x4_ASAP7_75t_R

MACRO AND2x6_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND2x6_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.554 0.243 ;
			RECT 0.31 0.027 0.554 0.045 ;
			RECT 0.45 0.027 0.468 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.028 0.252 0.15 ;
			RECT 0.072 0.028 0.252 0.046 ;
			RECT 0.072 0.028 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.107 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.231 0.243 ;
			RECT 0.18 0.064 0.198 0.243 ;
			RECT 0.179 0.182 0.306 0.2 ;
			RECT 0.288 0.121 0.306 0.2 ;
			RECT 0.115 0.064 0.198 0.082 ;

	END

END AND2x6_ASAP7_75t_R

MACRO AND3x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND3x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.183 0.306 0.201 ;
			RECT 0.288 0.076 0.306 0.201 ;
			RECT 0.261 0.076 0.306 0.094 ;
			RECT 0.261 0.183 0.279 0.235 ;
			RECT 0.261 0.034 0.279 0.094 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.263 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END AND3x1_ASAP7_75t_R

MACRO AND3x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND3x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.261 0.027 0.36 0.045 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END AND3x2_ASAP7_75t_R

MACRO AND3x4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND3x4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.23 0.243 ;
			RECT 0.018 0.027 0.23 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.189 0.649 0.207 ;
			RECT 0.612 0.099 0.649 0.117 ;
			RECT 0.612 0.099 0.63 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.189 0.541 0.207 ;
			RECT 0.504 0.099 0.541 0.117 ;
			RECT 0.504 0.099 0.522 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.26 0.225 0.746 0.243 ;
			RECT 0.728 0.027 0.746 0.243 ;
			RECT 0.26 0.042 0.278 0.243 ;
			RECT 0.218 0.126 0.278 0.144 ;
			RECT 0.634 0.027 0.746 0.045 ;
			RECT 0.472 0.063 0.701 0.081 ;
			RECT 0.31 0.027 0.554 0.045 ;

	END

END AND3x4_ASAP7_75t_R

MACRO AND4x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND4x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.299 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.164 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.234 0.189 0.306 0.207 ;
			RECT 0.288 0.12 0.306 0.207 ;
			RECT 0.018 0.027 0.085 0.045 ;

	END

END AND4x1_ASAP7_75t_R

MACRO AND4x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND4x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.164 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.153 0.189 0.171 0.243 ;
			RECT 0.099 0.189 0.171 0.207 ;
			RECT 0.099 0.119 0.117 0.207 ;
			RECT 0.364 0.027 0.414 0.045 ;

	END

END AND4x2_ASAP7_75t_R

MACRO AND5x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND5x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.349 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.35 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.164 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.288 0.189 0.36 0.207 ;
			RECT 0.342 0.116 0.36 0.207 ;
			RECT 0.018 0.027 0.07 0.045 ;

	END

END AND5x1_ASAP7_75t_R

MACRO AND5x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AND5x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.958 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.958 0.027 1.062 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.72 0.189 0.757 0.207 ;
			RECT 0.72 0.099 0.757 0.117 ;
			RECT 0.72 0.099 0.738 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.593 0.189 0.63 0.207 ;
			RECT 0.612 0.099 0.63 0.207 ;
			RECT 0.593 0.099 0.63 0.117 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.189 0.487 0.207 ;
			RECT 0.45 0.099 0.487 0.117 ;
			RECT 0.45 0.099 0.468 0.207 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.269 0.189 0.306 0.207 ;
			RECT 0.288 0.099 0.306 0.207 ;
			RECT 0.269 0.099 0.306 0.117 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.225 0.9 0.243 ;
			RECT 0.882 0.027 0.9 0.243 ;
			RECT 0.882 0.126 0.942 0.144 ;
			RECT 0.742 0.027 0.9 0.045 ;
			RECT 0.58 0.063 0.824 0.081 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.256 0.063 0.5 0.081 ;
			RECT 0.094 0.027 0.338 0.045 ;

	END

END AND5x2_ASAP7_75t_R

MACRO AO211x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO211x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.742 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.311 0.144 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.215 0.063 0.252 0.081 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.153 0.541 0.171 ;
			RECT 0.504 0.063 0.522 0.171 ;
			RECT 0.485 0.063 0.522 0.081 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.666 0.125 0.743 0.143 ;
			RECT 0.094 0.027 0.684 0.045 ;
			RECT 0.31 0.189 0.608 0.207 ;
			RECT 0.04 0.225 0.393 0.243 ;

	END

END AO211x2_ASAP7_75t_R

MACRO AO21x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO21x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.23 0.225 0.295 0.243 ;
			RECT 0.277 0.038 0.295 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.189 0.252 0.207 ;
			RECT 0.234 0.027 0.252 0.207 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AO21x1_ASAP7_75t_R

MACRO AO21x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO21x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.23 0.225 0.333 0.243 ;
			RECT 0.315 0.069 0.333 0.243 ;
			RECT 0.276 0.069 0.333 0.087 ;
			RECT 0.276 0.038 0.294 0.087 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.189 0.252 0.207 ;
			RECT 0.234 0.027 0.252 0.207 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AO21x2_ASAP7_75t_R

MACRO AO221x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO221x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.459 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.126 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;
			RECT 0.396 0.126 0.474 0.144 ;
			RECT 0.396 0.027 0.414 0.144 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.2 0.189 0.339 0.207 ;
			RECT 0.039 0.225 0.176 0.243 ;

	END

END AO221x1_ASAP7_75t_R

MACRO AO221x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO221x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.549 0.243 ;
			RECT 0.531 0.027 0.549 0.243 ;
			RECT 0.459 0.027 0.549 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.126 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;
			RECT 0.396 0.126 0.474 0.144 ;
			RECT 0.396 0.027 0.414 0.144 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.2 0.189 0.339 0.207 ;
			RECT 0.039 0.225 0.176 0.243 ;

	END

END AO221x2_ASAP7_75t_R

MACRO AO222x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO222x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.526 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.531 0.027 0.63 0.045 ;
			RECT 0.531 0.027 0.549 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.009 0.189 0.122 0.207 ;
			RECT 0.009 0.027 0.027 0.207 ;
			RECT 0.486 0.126 0.554 0.144 ;
			RECT 0.486 0.027 0.504 0.144 ;
			RECT 0.009 0.027 0.504 0.045 ;
			RECT 0.342 0.225 0.468 0.243 ;
			RECT 0.342 0.189 0.36 0.243 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO222x2_ASAP7_75t_R

MACRO AO22x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO22x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.418 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.287 0.081 ;
			RECT 0.234 0.063 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.342 0.126 0.419 0.144 ;
			RECT 0.107 0.027 0.36 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO22x1_ASAP7_75t_R

MACRO AO22x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO22x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.418 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.287 0.081 ;
			RECT 0.234 0.063 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.342 0.126 0.419 0.144 ;
			RECT 0.107 0.027 0.36 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO22x2_ASAP7_75t_R

MACRO AO31x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO31x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.741 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.742 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.099 0.576 0.149 ;
			RECT 0.504 0.099 0.576 0.117 ;
			RECT 0.485 0.153 0.522 0.171 ;
			RECT 0.504 0.099 0.522 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.414 0.149 ;
			RECT 0.288 0.099 0.414 0.117 ;
			RECT 0.288 0.153 0.325 0.171 ;
			RECT 0.288 0.07 0.306 0.171 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.059 0.207 ;
			RECT 0.018 0.027 0.059 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.612 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.612 0.189 0.63 0.243 ;
			RECT 0.199 0.189 0.63 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.666 0.126 0.797 0.144 ;
			RECT 0.2 0.063 0.252 0.081 ;
			RECT 0.526 0.027 0.684 0.045 ;
			RECT 0.364 0.063 0.608 0.081 ;
			RECT 0.04 0.225 0.554 0.243 ;
			RECT 0.094 0.027 0.447 0.045 ;

	END

END AO31x2_ASAP7_75t_R

MACRO AO322x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO322x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.634 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.634 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.153 0.325 0.171 ;
			RECT 0.288 0.063 0.325 0.081 ;
			RECT 0.288 0.063 0.306 0.171 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.063 0.541 0.081 ;
			RECT 0.504 0.063 0.522 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.396 0.189 0.576 0.207 ;
			RECT 0.558 0.126 0.576 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.558 0.126 0.743 0.144 ;
			RECT 0.04 0.027 0.446 0.045 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.189 0.198 0.243 ;
			RECT 0.18 0.189 0.338 0.207 ;
			RECT 0.256 0.225 0.5 0.243 ;

	END

END AO322x2_ASAP7_75t_R

MACRO AO32x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO32x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.063 0.063 0.081 ;
			RECT 0.045 0.034 0.063 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.062 0.126 0.108 0.144 ;
			RECT 0.09 0.027 0.108 0.144 ;
			RECT 0.09 0.027 0.414 0.045 ;
			RECT 0.148 0.225 0.392 0.243 ;

	END

END AO32x1_ASAP7_75t_R

MACRO AO32x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO32x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.068 0.117 0.086 ;
			RECT 0.099 0.037 0.117 0.086 ;
			RECT 0.018 0.068 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.189 0.33 0.207 ;
			RECT 0.288 0.07 0.306 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.364 0.189 0.468 0.207 ;
			RECT 0.45 0.027 0.468 0.207 ;
			RECT 0.093 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.468 0.045 ;
			RECT 0.202 0.225 0.446 0.243 ;

	END

END AO32x2_ASAP7_75t_R

MACRO AO331x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO331x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.081 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B3
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.072 0.063 0.09 0.152 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.522 0.045 ;
			RECT 0.308 0.189 0.447 0.207 ;
			RECT 0.146 0.225 0.393 0.243 ;

	END

END AO331x1_ASAP7_75t_R

MACRO AO331x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO331x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.027 0.135 0.045 ;
			RECT 0.072 0.225 0.122 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.126 0.063 0.144 0.152 ;
			RECT 0.126 0.063 0.198 0.081 ;
			RECT 0.18 0.027 0.198 0.081 ;
			RECT 0.18 0.027 0.576 0.045 ;
			RECT 0.362 0.189 0.501 0.207 ;
			RECT 0.2 0.225 0.447 0.243 ;

	END

END AO331x2_ASAP7_75t_R

MACRO AO332x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO332x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.094 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.072 0.063 0.09 0.151 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.576 0.045 ;
			RECT 0.146 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.234 0.189 0.393 0.207 ;
			RECT 0.308 0.225 0.556 0.243 ;

	END

END AO332x1_ASAP7_75t_R

MACRO AO332x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO332x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.148 0.045 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.189 0.63 0.207 ;
			RECT 0.612 0.027 0.63 0.207 ;
			RECT 0.126 0.063 0.144 0.151 ;
			RECT 0.126 0.063 0.198 0.081 ;
			RECT 0.18 0.027 0.198 0.081 ;
			RECT 0.18 0.027 0.63 0.045 ;
			RECT 0.2 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.288 0.189 0.447 0.207 ;
			RECT 0.362 0.225 0.61 0.243 ;

	END

END AO332x2_ASAP7_75t_R

MACRO AO333x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO333x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.081 0.045 ;
			RECT 0.018 0.225 0.069 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.063 0.09 0.152 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.63 0.045 ;
			RECT 0.31 0.189 0.576 0.207 ;
			RECT 0.148 0.225 0.395 0.243 ;

	END

END AO333x1_ASAP7_75t_R

MACRO AO333x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO333x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.081 0.117 0.099 ;
			RECT 0.099 0.045 0.117 0.099 ;
			RECT 0.018 0.081 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.07 0.63 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.067 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.684 0.045 ;
			RECT 0.364 0.189 0.63 0.207 ;
			RECT 0.202 0.225 0.449 0.243 ;

	END

END AO333x2_ASAP7_75t_R

MACRO AO33x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AO33x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.068 0.117 0.086 ;
			RECT 0.099 0.037 0.117 0.086 ;
			RECT 0.018 0.068 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.361 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.067 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.522 0.045 ;
			RECT 0.199 0.225 0.449 0.243 ;

	END

END AO33x2_ASAP7_75t_R

MACRO AOI211x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI211x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.519 0.189 0.63 0.207 ;
			RECT 0.612 0.027 0.63 0.207 ;
			RECT 0.091 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.126 0.229 0.144 ;
			RECT 0.18 0.189 0.223 0.207 ;
			RECT 0.18 0.063 0.22 0.081 ;
			RECT 0.18 0.063 0.198 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.123 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.153 0.442 0.171 ;
			RECT 0.396 0.063 0.442 0.081 ;
			RECT 0.396 0.063 0.414 0.171 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.126 0.554 0.144 ;
			RECT 0.504 0.063 0.55 0.081 ;
			RECT 0.504 0.063 0.522 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.288 0.189 0.449 0.207 ;
			RECT 0.361 0.225 0.608 0.243 ;

	END

END AOI211x1_ASAP7_75t_R

MACRO AOI211xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI211xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.04 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AOI211xp5_ASAP7_75t_R

MACRO AOI21x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI21x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.369 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.018 0.225 0.063 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.063 0.306 0.164 ;
			RECT 0.126 0.063 0.306 0.081 ;
			RECT 0.126 0.063 0.144 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.19 0.125 0.256 0.143 ;
			RECT 0.19 0.099 0.227 0.171 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.189 0.36 0.207 ;
			RECT 0.342 0.116 0.36 0.207 ;
			RECT 0.072 0.07 0.09 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.333 0.243 ;

	END

END AOI21x1_ASAP7_75t_R

MACRO AOI21xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI21xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.107 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END AOI21xp33_ASAP7_75t_R

MACRO AOI21xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI21xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.142 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.034 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END AOI21xp5_ASAP7_75t_R

MACRO AOI221x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI221x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.634 0.189 0.738 0.207 ;
			RECT 0.72 0.045 0.738 0.207 ;
			RECT 0.256 0.045 0.738 0.063 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.153 0.217 0.171 ;
			RECT 0.18 0.027 0.198 0.171 ;
			RECT 0.161 0.027 0.198 0.045 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.126 0.149 0.144 ;
			RECT 0.053 0.153 0.09 0.171 ;
			RECT 0.072 0.027 0.09 0.171 ;
			RECT 0.053 0.027 0.09 0.045 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.081 0.325 0.099 ;
			RECT 0.269 0.153 0.306 0.171 ;
			RECT 0.288 0.081 0.306 0.171 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.153 0.487 0.171 ;
			RECT 0.45 0.081 0.468 0.171 ;
			RECT 0.391 0.126 0.468 0.144 ;
			RECT 0.431 0.081 0.468 0.099 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.126 0.636 0.144 ;
			RECT 0.539 0.189 0.576 0.207 ;
			RECT 0.558 0.081 0.576 0.207 ;
			RECT 0.539 0.081 0.576 0.099 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.225 0.716 0.243 ;
			RECT 0.04 0.189 0.5 0.207 ;

	END

END AOI221x1_ASAP7_75t_R

MACRO AOI221xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI221xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.23 0.045 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.201 0.189 0.339 0.207 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AOI221xp5_ASAP7_75t_R

MACRO AOI222xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI222xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.399 0.045 ;
			RECT 0.018 0.189 0.122 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.034 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.342 0.225 0.468 0.243 ;
			RECT 0.342 0.189 0.36 0.243 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI222xp33_ASAP7_75t_R

MACRO AOI22x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI22x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.309 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.038 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.153 0.379 0.171 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.431 0.153 0.468 0.171 ;
			RECT 0.45 0.063 0.468 0.171 ;
			RECT 0.288 0.063 0.468 0.081 ;
			RECT 0.288 0.063 0.306 0.152 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.161 0.189 0.198 0.207 ;
			RECT 0.18 0.099 0.198 0.207 ;
			RECT 0.161 0.099 0.198 0.117 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.252 0.154 ;
			RECT 0.072 0.063 0.252 0.081 ;
			RECT 0.072 0.189 0.109 0.207 ;
			RECT 0.072 0.063 0.09 0.207 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.5 0.243 ;

	END

END AOI22x1_ASAP7_75t_R

MACRO AOI22xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI22xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI22xp33_ASAP7_75t_R

MACRO AOI22xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI22xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.07 0.144 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI22xp5_ASAP7_75t_R

MACRO AOI311xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI311xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.198 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.234 0.243 ;

	END

END AOI311xp33_ASAP7_75t_R

MACRO AOI31xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI31xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.201 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.093 0.225 0.23 0.243 ;

	END

END AOI31xp33_ASAP7_75t_R

MACRO AOI31xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI31xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.585 0.225 0.663 0.243 ;
			RECT 0.585 0.189 0.603 0.243 ;
			RECT 0.202 0.189 0.603 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.202 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.666 0.07 0.684 0.2 ;
			RECT 0.553 0.126 0.684 0.144 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.126 0.419 0.144 ;
			RECT 0.288 0.063 0.325 0.081 ;
			RECT 0.288 0.063 0.306 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.059 0.207 ;
			RECT 0.018 0.027 0.059 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.027 0.663 0.045 ;
			RECT 0.364 0.081 0.608 0.099 ;
			RECT 0.04 0.225 0.554 0.243 ;
			RECT 0.094 0.027 0.447 0.045 ;

	END

END AOI31xp67_ASAP7_75t_R

MACRO AOI321xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI321xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.198 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.225 0.396 0.243 ;
			RECT 0.094 0.189 0.23 0.207 ;

	END

END AOI321xp33_ASAP7_75t_R

MACRO AOI322xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI322xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.189 0.468 0.207 ;
			RECT 0.45 0.027 0.468 0.207 ;
			RECT 0.147 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.165 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.165 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.225 0.45 0.243 ;
			RECT 0.039 0.189 0.284 0.207 ;

	END

END AOI322xp5_ASAP7_75t_R

MACRO AOI32xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI32xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.04 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.058 0.243 ;
			RECT 0.018 0.063 0.058 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.104 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.104 0.063 0.144 0.081 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.222 0.207 ;
			RECT 0.18 0.07 0.198 0.207 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END AOI32xp33_ASAP7_75t_R

MACRO AOI331xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI331xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.417 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.201 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.189 0.393 0.207 ;
			RECT 0.092 0.225 0.339 0.243 ;

	END

END AOI331xp33_ASAP7_75t_R

MACRO AOI332xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI332xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.417 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.201 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.225 0.502 0.243 ;
			RECT 0.092 0.189 0.339 0.207 ;

	END

END AOI332xp33_ASAP7_75t_R

MACRO AOI333xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI333xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.413 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.201 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.225 0.515 0.243 ;
			RECT 0.094 0.189 0.34 0.207 ;

	END

END AOI333xp33_ASAP7_75t_R

MACRO AOI33xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN AOI33xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.201 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.338 0.243 ;

	END

END AOI33xp33_ASAP7_75t_R

MACRO BUFx10_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx10_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.199 0.027 0.738 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.689 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx10_ASAP7_75t_R

MACRO BUFx12_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx12_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.199 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.8 0.144 ;
			RECT 0.094 0.027 0.144 0.045 ;

	END

END BUFx12_ASAP7_75t_R

MACRO BUFx12f_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx12f_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.972 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.31 0.027 0.954 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.074 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.972 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.972 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.243 ;
			RECT 0.261 0.126 0.311 0.144 ;
			RECT 0.094 0.027 0.279 0.045 ;

	END

END BUFx12f_ASAP7_75t_R

MACRO BUFx16f_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx16f_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 1.17 0.243 ;
			RECT 1.152 0.027 1.17 0.243 ;
			RECT 0.31 0.027 1.17 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.06 0.243 ;
			RECT 0.018 0.027 0.06 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.234 0.126 1.124 0.144 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END BUFx16f_ASAP7_75t_R

MACRO BUFx24_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx24_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.62 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 1.602 0.243 ;
			RECT 1.584 0.027 1.602 0.243 ;
			RECT 0.31 0.027 1.602 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.62 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.62 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.234 0.126 1.553 0.144 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END BUFx24_ASAP7_75t_R

MACRO BUFx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.145 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.203 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx2_ASAP7_75t_R

MACRO BUFx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.145 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.26 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx3_ASAP7_75t_R

MACRO BUFx4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.357 0.243 ;
			RECT 0.339 0.027 0.357 0.243 ;
			RECT 0.145 0.027 0.357 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.314 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx4_ASAP7_75t_R

MACRO BUFx4f_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx4f_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.199 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.098 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.367 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx4f_ASAP7_75t_R

MACRO BUFx5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.145 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.368 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx5_ASAP7_75t_R

MACRO BUFx6f_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx6f_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.202 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.473 0.144 ;
			RECT 0.094 0.027 0.144 0.045 ;

	END

END BUFx6f_ASAP7_75t_R

MACRO BUFx8_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN BUFx8_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.202 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.098 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.581 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx8_ASAP7_75t_R

MACRO CKINVDCx10_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx10_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.296 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.224 0.243 ;
			RECT 1.206 0.063 1.224 0.243 ;
			RECT 1.174 0.063 1.224 0.081 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.17 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.296 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.296 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx10_ASAP7_75t_R

MACRO CKINVDCx11_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx11_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.31 0.243 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.354 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx11_ASAP7_75t_R

MACRO CKINVDCx12_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx12_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.31 0.243 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.354 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx12_ASAP7_75t_R

MACRO CKINVDCx14_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx14_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.512 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.44 0.243 ;
			RECT 1.422 0.063 1.44 0.243 ;
			RECT 1.39 0.063 1.44 0.081 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.397 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.512 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.512 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx14_ASAP7_75t_R

MACRO CKINVDCx16_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx16_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.62 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 1.548 0.243 ;
			RECT 1.53 0.063 1.548 0.243 ;
			RECT 1.498 0.063 1.548 0.081 ;
			RECT 1.368 0.063 1.418 0.081 ;
			RECT 1.368 0.063 1.386 0.243 ;
			RECT 1.098 0.063 1.116 0.243 ;
			RECT 1.066 0.063 1.116 0.081 ;
			RECT 0.936 0.063 0.986 0.081 ;
			RECT 0.936 0.063 0.954 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.634 0.063 0.684 0.081 ;
			RECT 0.504 0.063 0.554 0.081 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.202 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.122 0.081 ;
			RECT 0.072 0.063 0.09 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.412 0.126 1.505 0.144 ;
			RECT 1.444 0.027 1.462 0.144 ;
			RECT 0.158 0.027 1.462 0.045 ;
			RECT 0.98 0.126 1.072 0.144 ;
			RECT 1.017 0.027 1.035 0.144 ;
			RECT 0.547 0.126 0.639 0.144 ;
			RECT 0.584 0.027 0.602 0.144 ;
			RECT 0.126 0.126 0.208 0.144 ;
			RECT 0.158 0.027 0.176 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.62 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.62 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.26 0.126 1.316 0.144 ;
			RECT 1.26 0.09 1.278 0.144 ;
			RECT 1.174 0.09 1.326 0.108 ;
			RECT 1.155 0.162 1.31 0.18 ;
			RECT 1.206 0.126 1.224 0.18 ;
			RECT 1.166 0.126 1.224 0.144 ;
			RECT 0.742 0.162 0.897 0.18 ;
			RECT 0.828 0.126 0.846 0.18 ;
			RECT 0.828 0.126 0.886 0.144 ;
			RECT 0.736 0.126 0.792 0.144 ;
			RECT 0.774 0.09 0.792 0.144 ;
			RECT 0.726 0.09 0.878 0.108 ;
			RECT 0.31 0.162 0.465 0.18 ;
			RECT 0.396 0.126 0.414 0.18 ;
			RECT 0.396 0.126 0.454 0.144 ;
			RECT 0.304 0.126 0.36 0.144 ;
			RECT 0.342 0.09 0.36 0.144 ;
			RECT 0.294 0.09 0.446 0.108 ;

	END

END CKINVDCx16_ASAP7_75t_R

MACRO CKINVDCx20_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx20_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.052 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 1.98 0.243 ;
			RECT 1.962 0.063 1.98 0.243 ;
			RECT 1.93 0.063 1.98 0.081 ;
			RECT 1.8 0.063 1.85 0.081 ;
			RECT 1.8 0.063 1.818 0.243 ;
			RECT 1.53 0.063 1.548 0.243 ;
			RECT 1.498 0.063 1.548 0.081 ;
			RECT 1.368 0.063 1.418 0.081 ;
			RECT 1.368 0.063 1.386 0.243 ;
			RECT 1.098 0.063 1.116 0.243 ;
			RECT 1.066 0.063 1.116 0.081 ;
			RECT 0.936 0.063 0.986 0.081 ;
			RECT 0.936 0.063 0.954 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.634 0.063 0.684 0.081 ;
			RECT 0.504 0.063 0.554 0.081 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.202 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.122 0.081 ;
			RECT 0.072 0.063 0.09 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.844 0.126 1.937 0.144 ;
			RECT 1.876 0.027 1.894 0.144 ;
			RECT 0.158 0.027 1.894 0.045 ;
			RECT 1.412 0.126 1.505 0.144 ;
			RECT 1.444 0.027 1.462 0.144 ;
			RECT 0.98 0.126 1.072 0.144 ;
			RECT 1.017 0.027 1.035 0.144 ;
			RECT 0.547 0.126 0.639 0.144 ;
			RECT 0.584 0.027 0.602 0.144 ;
			RECT 0.126 0.126 0.208 0.144 ;
			RECT 0.158 0.027 0.176 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.052 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.052 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.692 0.126 1.748 0.144 ;
			RECT 1.692 0.09 1.71 0.144 ;
			RECT 1.606 0.09 1.758 0.108 ;
			RECT 1.587 0.162 1.742 0.18 ;
			RECT 1.638 0.126 1.656 0.18 ;
			RECT 1.598 0.126 1.656 0.144 ;
			RECT 1.26 0.126 1.316 0.144 ;
			RECT 1.26 0.09 1.278 0.144 ;
			RECT 1.174 0.09 1.326 0.108 ;
			RECT 1.155 0.162 1.31 0.18 ;
			RECT 1.206 0.126 1.224 0.18 ;
			RECT 1.166 0.126 1.224 0.144 ;
			RECT 0.742 0.162 0.897 0.18 ;
			RECT 0.828 0.126 0.846 0.18 ;
			RECT 0.828 0.126 0.886 0.144 ;
			RECT 0.736 0.126 0.792 0.144 ;
			RECT 0.774 0.09 0.792 0.144 ;
			RECT 0.726 0.09 0.878 0.108 ;
			RECT 0.31 0.162 0.465 0.18 ;
			RECT 0.396 0.126 0.414 0.18 ;
			RECT 0.396 0.126 0.454 0.144 ;
			RECT 0.304 0.126 0.36 0.144 ;
			RECT 0.342 0.09 0.36 0.144 ;
			RECT 0.294 0.09 0.446 0.108 ;

	END

END CKINVDCx20_ASAP7_75t_R

MACRO CKINVDCx5p33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx5p33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.094 0.243 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.138 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx5p33_ASAP7_75t_R

MACRO CKINVDCx6p67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx6p67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.296 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.224 0.243 ;
			RECT 1.206 0.063 1.224 0.243 ;
			RECT 1.174 0.063 1.224 0.081 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.17 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.296 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.296 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx6p67_ASAP7_75t_R

MACRO CKINVDCx8_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx8_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.094 0.243 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.138 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx8_ASAP7_75t_R

MACRO CKINVDCx9p33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN CKINVDCx9p33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.512 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.44 0.243 ;
			RECT 1.422 0.063 1.44 0.243 ;
			RECT 1.39 0.063 1.44 0.081 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.397 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.512 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.512 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx9p33_ASAP7_75t_R

MACRO DECAPx10_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN DECAPx10_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.558 0.045 0.576 0.15 ;
			RECT 0.558 0.045 1.148 0.063 ;
			RECT 0.04 0.207 0.63 0.225 ;
			RECT 0.612 0.121 0.63 0.225 ;

	END

END DECAPx10_ASAP7_75t_R

MACRO DECAPx1_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN DECAPx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.207 0.144 0.225 ;
			RECT 0.126 0.121 0.144 0.225 ;
			RECT 0.072 0.045 0.09 0.15 ;
			RECT 0.072 0.045 0.122 0.063 ;

	END

END DECAPx1_ASAP7_75t_R

MACRO DECAPx2_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN DECAPx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.045 0.144 0.15 ;
			RECT 0.126 0.045 0.284 0.063 ;
			RECT 0.04 0.207 0.198 0.225 ;
			RECT 0.18 0.121 0.198 0.225 ;

	END

END DECAPx2_ASAP7_75t_R

MACRO DECAPx2b_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN DECAPx2b_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.162 0.249 0.18 ;
			RECT 0.18 0.126 0.198 0.18 ;
			RECT 0.18 0.126 0.238 0.144 ;
			RECT 0.088 0.126 0.144 0.144 ;
			RECT 0.126 0.09 0.144 0.144 ;
			RECT 0.078 0.09 0.23 0.108 ;

	END

END DECAPx2b_ASAP7_75t_R

MACRO DECAPx4_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN DECAPx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.234 0.045 0.252 0.15 ;
			RECT 0.234 0.045 0.5 0.063 ;
			RECT 0.04 0.207 0.306 0.225 ;
			RECT 0.288 0.121 0.306 0.225 ;

	END

END DECAPx4_ASAP7_75t_R

MACRO DECAPx6_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN DECAPx6_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.342 0.045 0.36 0.15 ;
			RECT 0.342 0.045 0.716 0.063 ;
			RECT 0.04 0.207 0.414 0.225 ;
			RECT 0.396 0.121 0.414 0.225 ;

	END

END DECAPx6_ASAP7_75t_R

MACRO DFFASRHQNx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFASRHQNx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.336 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.336 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.182 0.117 0.236 ;
			RECT 0.072 0.182 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN RESETN
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.632 0.144 1.067 0.162 ;
			LAYER M1 ;
			RECT 1.044 0.102 1.062 0.167 ;
			RECT 0.612 0.072 0.668 0.09 ;
			RECT 0.612 0.144 0.662 0.162 ;
			RECT 0.612 0.072 0.63 0.162 ;
			LAYER V1 ;
			RECT 0.637 0.144 0.655 0.162 ;
			RECT 1.044 0.144 1.062 0.162 ;

		END 

	END RESETN
	PIN SETN
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.783 0.18 1.067 0.198 ;
			LAYER M1 ;
			RECT 0.774 0.18 0.811 0.198 ;
			RECT 0.774 0.097 0.792 0.198 ;
			LAYER V1 ;
			RECT 0.788 0.18 0.806 0.198 ;

		END 

	END SETN
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.963 0.036 0.981 0.234 ;
			RECT 0.963 0.036 1.008 0.054 ;
			RECT 0.855 0.222 0.936 0.24 ;
			RECT 0.918 0.053 0.936 0.24 ;
			RECT 0.693 0.036 0.711 0.212 ;
			RECT 0.558 0.036 0.576 0.106 ;
			RECT 0.558 0.036 0.77 0.054 ;
			RECT 0.486 0.18 0.547 0.198 ;
			RECT 0.486 0.027 0.504 0.198 ;
			RECT 0.418 0.027 0.504 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.142 0.027 0.198 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.018 0.108 0.047 0.126 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 1.314 0.103 1.332 0.18 ;
			RECT 1.17 0.216 1.202 0.234 ;
			RECT 1.098 0.102 1.116 0.167 ;
			RECT 0.882 0.067 0.9 0.173 ;
			RECT 0.829 0.103 0.847 0.171 ;
			RECT 0.778 0.216 0.819 0.234 ;
			RECT 0.729 0.137 0.747 0.203 ;
			RECT 0.415 0.225 0.608 0.243 ;
			RECT 0.45 0.103 0.468 0.151 ;
			RECT 0.396 0.067 0.414 0.15 ;
			RECT 0.369 0.169 0.387 0.216 ;
			RECT 0.342 0.103 0.36 0.15 ;
			RECT 0.142 0.07 0.16 0.164 ;
			LAYER M2 ;
			RECT 0.913 0.108 1.337 0.126 ;
			RECT 0.783 0.216 1.198 0.234 ;
			RECT 0.741 0.036 1.008 0.054 ;
			RECT 0.018 0.072 0.926 0.09 ;
			RECT 0.175 0.108 0.852 0.126 ;
			RECT 0.364 0.18 0.752 0.198 ;
			LAYER V1 ;
			RECT 1.314 0.108 1.332 0.126 ;
			RECT 1.175 0.216 1.193 0.234 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 0.985 0.036 1.003 0.054 ;
			RECT 0.918 0.108 0.936 0.126 ;
			RECT 0.882 0.072 0.9 0.09 ;
			RECT 0.829 0.108 0.847 0.126 ;
			RECT 0.788 0.216 0.806 0.234 ;
			RECT 0.746 0.036 0.764 0.054 ;
			RECT 0.729 0.18 0.747 0.198 ;
			RECT 0.512 0.18 0.53 0.198 ;
			RECT 0.45 0.108 0.468 0.126 ;
			RECT 0.396 0.072 0.414 0.09 ;
			RECT 0.369 0.18 0.387 0.198 ;
			RECT 0.342 0.108 0.36 0.126 ;
			RECT 0.18 0.108 0.198 0.126 ;
			RECT 0.142 0.072 0.16 0.09 ;
			RECT 0.018 0.072 0.036 0.09 ;

	END

END DFFASRHQNx1_ASAP7_75t_R

MACRO DFFHQNx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFHQNx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 1.012 0.027 1.062 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx1_ASAP7_75t_R

MACRO DFFHQNx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFHQNx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.216 1.117 0.234 ;
			RECT 1.099 0.036 1.117 0.234 ;
			RECT 1.012 0.036 1.117 0.054 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx2_ASAP7_75t_R

MACRO DFFHQNx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFHQNx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.171 0.243 ;
			RECT 1.153 0.027 1.171 0.243 ;
			RECT 1.012 0.027 1.171 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx3_ASAP7_75t_R

MACRO DFFHQx4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFHQx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.125 0.225 1.333 0.243 ;
			RECT 1.313 0.027 1.333 0.243 ;
			RECT 1.125 0.027 1.333 0.045 ;
			RECT 1.125 0.201 1.143 0.243 ;
			RECT 1.125 0.027 1.143 0.069 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.012 0.225 1.098 0.243 ;
			RECT 1.08 0.027 1.098 0.243 ;
			RECT 1.08 0.127 1.175 0.145 ;
			RECT 1.012 0.027 1.098 0.045 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQx4_ASAP7_75t_R

MACRO DFFLQNx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFLQNx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 1.012 0.027 1.062 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx1_ASAP7_75t_R

MACRO DFFLQNx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFLQNx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.115 0.243 ;
			RECT 1.097 0.027 1.115 0.243 ;
			RECT 1.012 0.027 1.115 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx2_ASAP7_75t_R

MACRO DFFLQNx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFLQNx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.171 0.243 ;
			RECT 1.153 0.027 1.171 0.243 ;
			RECT 1.011 0.027 1.171 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx3_ASAP7_75t_R

MACRO DFFLQx4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DFFLQx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.125 0.225 1.333 0.243 ;
			RECT 1.313 0.027 1.333 0.243 ;
			RECT 1.125 0.027 1.333 0.045 ;
			RECT 1.125 0.201 1.143 0.243 ;
			RECT 1.125 0.027 1.143 0.069 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.012 0.225 1.098 0.243 ;
			RECT 1.08 0.027 1.098 0.243 ;
			RECT 1.08 0.127 1.175 0.145 ;
			RECT 1.012 0.027 1.098 0.045 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQx4_ASAP7_75t_R

MACRO DHLx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DHLx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.742 0.027 0.792 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.72 0.122 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.743 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx1_ASAP7_75t_R

MACRO DHLx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DHLx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.741 0.216 0.85 0.234 ;
			RECT 0.832 0.036 0.85 0.234 ;
			RECT 0.742 0.036 0.85 0.054 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.72 0.09 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.797 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx2_ASAP7_75t_R

MACRO DHLx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DHLx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.918 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.688 0.225 0.9 0.243 ;
			RECT 0.882 0.027 0.9 0.243 ;
			RECT 0.688 0.027 0.9 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.918 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.918 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.828 0.09 0.846 0.167 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.72 0.09 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.851 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx3_ASAP7_75t_R

MACRO DLLx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DLLx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.735 0.027 0.792 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.72 0.106 0.738 0.2 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.743 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx1_ASAP7_75t_R

MACRO DLLx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DLLx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.688 0.225 0.847 0.243 ;
			RECT 0.829 0.027 0.847 0.243 ;
			RECT 0.688 0.027 0.847 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.8 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx2_ASAP7_75t_R

MACRO DLLx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN DLLx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.918 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.216 0.901 0.234 ;
			RECT 0.882 0.036 0.901 0.234 ;
			RECT 0.742 0.036 0.901 0.054 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.918 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.918 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.8 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx3_ASAP7_75t_R

MACRO FAx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN FAx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN CON
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.128 0.072 0.543 0.09 ;
			LAYER M1 ;
			RECT 0.515 0.072 0.543 0.09 ;
			RECT 0.504 0.09 0.533 0.108 ;
			RECT 0.504 0.09 0.522 0.149 ;
			RECT 0.124 0.072 0.282 0.09 ;
			RECT 0.124 0.189 0.23 0.207 ;
			RECT 0.124 0.072 0.142 0.207 ;
			LAYER V1 ;
			RECT 0.133 0.072 0.151 0.09 ;
			RECT 0.52 0.072 0.538 0.09 ;

		END 

	END CON
	PIN SN
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.324 0.225 0.495 0.243 ;
			RECT 0.477 0.184 0.495 0.243 ;
			RECT 0.477 0.027 0.495 0.068 ;
			RECT 0.324 0.027 0.495 0.045 ;
			RECT 0.324 0.027 0.342 0.243 ;

		END 

	END SN
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.059 0.18 0.627 0.198 ;
			LAYER M1 ;
			RECT 0.599 0.18 0.63 0.198 ;
			RECT 0.612 0.121 0.63 0.198 ;
			RECT 0.383 0.18 0.414 0.198 ;
			RECT 0.396 0.121 0.414 0.198 ;
			RECT 0.059 0.18 0.09 0.198 ;
			RECT 0.072 0.121 0.09 0.198 ;
			LAYER V1 ;
			RECT 0.064 0.18 0.082 0.198 ;
			RECT 0.388 0.18 0.406 0.198 ;
			RECT 0.604 0.18 0.622 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.167 0.144 0.689 0.162 ;
			LAYER M1 ;
			RECT 0.666 0.121 0.684 0.167 ;
			RECT 0.288 0.121 0.306 0.167 ;
			RECT 0.167 0.144 0.198 0.162 ;
			RECT 0.18 0.121 0.198 0.162 ;
			LAYER V1 ;
			RECT 0.172 0.144 0.19 0.162 ;
			RECT 0.288 0.144 0.306 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;

		END 

	END B
	PIN CI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.108 0.587 0.126 ;
			LAYER M1 ;
			RECT 0.558 0.108 0.587 0.126 ;
			RECT 0.558 0.108 0.576 0.149 ;
			RECT 0.45 0.103 0.468 0.149 ;
			RECT 0.226 0.108 0.263 0.126 ;
			RECT 0.234 0.108 0.252 0.149 ;
			LAYER V1 ;
			RECT 0.234 0.108 0.252 0.126 ;
			RECT 0.45 0.108 0.468 0.126 ;
			RECT 0.564 0.108 0.582 0.126 ;

		END 

	END CI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.027 0.662 0.045 ;
			RECT 0.526 0.225 0.662 0.243 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END FAx1_ASAP7_75t_R

MACRO FILLER_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN FILLER_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.108 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.108 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.108 0.279 ;

		END 

	END VDD

END FILLER_ASAP7_75t_R

MACRO FILLERxp5_ASAP7_75t_R
	CLASS CORE SPACER ;
	FOREIGN FILLERxp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.054 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.054 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.054 0.279 ;

		END 

	END VDD

END FILLERxp5_ASAP7_75t_R

MACRO HAxp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN HAxp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN CON
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.162 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.075 0.18 0.243 ;

		END 

	END CON
	PIN SN
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.423 0.027 0.468 0.045 ;

		END 

	END SN
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.15 ;
			RECT 0.207 0.063 0.36 0.081 ;
			RECT 0.207 0.027 0.225 0.081 ;
			RECT 0.018 0.027 0.225 0.045 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.027 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.106 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.387 0.045 ;

	END

END HAxp5_ASAP7_75t_R

MACRO HB1xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN HB1xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.117 0.243 ;
			RECT 0.099 0.153 0.117 0.243 ;
			RECT 0.099 0.153 0.144 0.171 ;
			RECT 0.126 0.099 0.144 0.171 ;
			RECT 0.099 0.099 0.144 0.117 ;
			RECT 0.099 0.027 0.117 0.117 ;
			RECT 0.04 0.027 0.117 0.045 ;

	END

END HB1xp67_ASAP7_75t_R

MACRO HB2xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN HB2xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.202 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.04 0.027 0.144 0.045 ;

	END

END HB2xp67_ASAP7_75t_R

MACRO HB3xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN HB3xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.256 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.18 0.126 0.257 0.144 ;
			RECT 0.04 0.027 0.198 0.045 ;

	END

END HB3xp67_ASAP7_75t_R

MACRO HB4xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN HB4xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.081 0.055 0.099 ;
			RECT 0.018 0.081 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.18 0.126 0.311 0.144 ;
			RECT 0.04 0.027 0.198 0.045 ;

	END

END HB4xp67_ASAP7_75t_R

MACRO ICGx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.972 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.879 0.027 0.954 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.972 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.972 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx1_ASAP7_75t_R

MACRO ICGx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.026 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 1.008 0.243 ;
			RECT 0.99 0.027 1.008 0.243 ;
			RECT 0.879 0.027 1.008 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.026 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.026 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx2_ASAP7_75t_R

MACRO ICGx2p67DC_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx2p67DC_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx2p67DC_ASAP7_75t_R

MACRO ICGx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.879 0.027 1.062 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx3_ASAP7_75t_R

MACRO ICGx4DC_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx4DC_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx4DC_ASAP7_75t_R

MACRO ICGx4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.89 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.889 0.027 1.062 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx4_ASAP7_75t_R

MACRO ICGx5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.89 0.225 1.17 0.243 ;
			RECT 1.152 0.027 1.17 0.243 ;
			RECT 0.889 0.027 1.17 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx5_ASAP7_75t_R

MACRO ICGx5p33DC_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx5p33DC_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx5p33DC_ASAP7_75t_R

MACRO ICGx6p67DC_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx6p67DC_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx6p67DC_ASAP7_75t_R

MACRO ICGx8DC_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN ICGx8DC_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx8DC_ASAP7_75t_R

MACRO INVx11_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx11_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.094 0.027 0.684 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD

END INVx11_ASAP7_75t_R

MACRO INVx13_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx13_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.094 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD

END INVx13_ASAP7_75t_R

MACRO INVx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVx1_ASAP7_75t_R

MACRO INVx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END INVx2_ASAP7_75t_R

MACRO INVx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.094 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END INVx3_ASAP7_75t_R

MACRO INVx4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END INVx4_ASAP7_75t_R

MACRO INVx5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.094 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END INVx5_ASAP7_75t_R

MACRO INVx6_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx6_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.094 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD

END INVx6_ASAP7_75t_R

MACRO INVx8_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVx8_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.094 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD

END INVx8_ASAP7_75t_R

MACRO INVxp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVxp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVxp33_ASAP7_75t_R

MACRO INVxp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN INVxp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVxp67_ASAP7_75t_R

MACRO MAJIxp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN MAJIxp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.255 0.189 0.361 0.207 ;
			RECT 0.343 0.063 0.361 0.207 ;
			RECT 0.255 0.063 0.361 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.126 0.257 0.144 ;
			RECT 0.018 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.027 0.338 0.045 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END MAJIxp5_ASAP7_75t_R

MACRO MAJx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN MAJx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.364 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.333 0.207 ;
			RECT 0.315 0.106 0.333 0.207 ;
			RECT 0.283 0.126 0.333 0.144 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.121 0.126 0.198 0.144 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.063 0.036 0.207 ;
			RECT 0.368 0.063 0.386 0.149 ;
			RECT 0.018 0.063 0.386 0.081 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END MAJx2_ASAP7_75t_R

MACRO MAJx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN MAJx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.504 0.243 ;
			RECT 0.364 0.027 0.504 0.045 ;
			RECT 0.45 0.027 0.468 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.333 0.207 ;
			RECT 0.315 0.106 0.333 0.207 ;
			RECT 0.283 0.126 0.333 0.144 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.121 0.126 0.198 0.144 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.063 0.036 0.207 ;
			RECT 0.368 0.063 0.386 0.149 ;
			RECT 0.018 0.063 0.386 0.081 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END MAJx3_ASAP7_75t_R

MACRO NAND2x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND2x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.202 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.065 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END NAND2x1_ASAP7_75t_R

MACRO NAND2x1p5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND2x1p5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.261 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.063 0.338 0.081 ;
			RECT 0.094 0.027 0.225 0.045 ;

	END

END NAND2x1p5_ASAP7_75t_R

MACRO NAND2x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND2x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.418 0.063 0.522 0.081 ;
			RECT 0.018 0.063 0.122 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.242 0.189 0.279 0.207 ;
			RECT 0.261 0.106 0.279 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.177 ;
			RECT 0.322 0.099 0.468 0.117 ;
			RECT 0.322 0.063 0.34 0.117 ;
			RECT 0.2 0.063 0.34 0.081 ;
			RECT 0.072 0.099 0.218 0.117 ;
			RECT 0.2 0.063 0.218 0.117 ;
			RECT 0.072 0.189 0.109 0.207 ;
			RECT 0.072 0.099 0.09 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.5 0.045 ;

	END

END NAND2x2_ASAP7_75t_R

MACRO NAND2xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND2xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.143 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NAND2xp33_ASAP7_75t_R

MACRO NAND2xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND2xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.143 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.106 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NAND2xp5_ASAP7_75t_R

MACRO NAND2xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND2xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.202 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.106 0.252 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END NAND2xp67_ASAP7_75t_R

MACRO NAND3x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND3x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.418 0.063 0.576 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.402 0.18 0.468 0.198 ;
			RECT 0.45 0.108 0.468 0.198 ;
			RECT 0.4 0.108 0.468 0.126 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.243 0.18 0.306 0.198 ;
			RECT 0.288 0.108 0.306 0.198 ;
			RECT 0.246 0.108 0.306 0.126 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.061 0.103 0.079 0.203 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.5 0.045 ;
			RECT 0.094 0.063 0.338 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END NAND3x1_ASAP7_75t_R

MACRO NAND3x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND3x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 1.062 0.243 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.904 0.063 1.062 0.081 ;
			RECT 0.018 0.063 0.176 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.169 0.18 0.908 0.198 ;
			LAYER M1 ;
			RECT 0.866 0.189 0.903 0.207 ;
			RECT 0.885 0.108 0.903 0.207 ;
			RECT 0.174 0.189 0.211 0.207 ;
			RECT 0.174 0.106 0.192 0.207 ;
			LAYER V1 ;
			RECT 0.174 0.18 0.192 0.198 ;
			RECT 0.885 0.18 0.903 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.338 0.189 0.743 0.207 ;
			RECT 0.725 0.106 0.743 0.207 ;
			RECT 0.338 0.106 0.356 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.547 0.106 0.565 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.742 0.027 0.986 0.045 ;
			RECT 0.256 0.063 0.824 0.081 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.094 0.027 0.338 0.045 ;

	END

END NAND3x2_ASAP7_75t_R

MACRO NAND3xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND3xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END NAND3xp33_ASAP7_75t_R

MACRO NAND4xp25_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND4xp25_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.256 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END NAND4xp25_ASAP7_75t_R

MACRO NAND4xp75_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND4xp75_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.738 0.243 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.58 0.063 0.738 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.106 0.63 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.101 0.549 0.119 ;
			RECT 0.531 0.07 0.549 0.119 ;
			RECT 0.504 0.101 0.522 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.101 0.306 0.2 ;
			RECT 0.207 0.101 0.306 0.119 ;
			RECT 0.207 0.07 0.225 0.119 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.057 0.243 ;
			RECT 0.018 0.027 0.057 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.412 0.027 0.666 0.045 ;
			RECT 0.256 0.063 0.499 0.081 ;
			RECT 0.092 0.027 0.34 0.045 ;

	END

END NAND4xp75_ASAP7_75t_R

MACRO NAND5xp2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NAND5xp2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.009 0.225 0.317 0.243 ;
			RECT 0.009 0.027 0.07 0.045 ;
			RECT 0.009 0.027 0.027 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.2 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END NAND5xp2_ASAP7_75t_R

MACRO NOR2x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR2x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.23 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END NOR2x1_ASAP7_75t_R

MACRO NOR2x1p5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR2x1p5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.094 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.063 0.163 0.081 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.338 0.207 ;
			RECT 0.094 0.225 0.225 0.243 ;

	END

END NOR2x1p5_ASAP7_75t_R

MACRO NOR2x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR2x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.018 0.027 0.522 0.045 ;
			RECT 0.018 0.189 0.122 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.063 0.279 0.164 ;
			RECT 0.242 0.063 0.279 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.322 0.153 0.468 0.171 ;
			RECT 0.45 0.093 0.468 0.171 ;
			RECT 0.2 0.189 0.34 0.207 ;
			RECT 0.322 0.153 0.34 0.207 ;
			RECT 0.2 0.153 0.218 0.207 ;
			RECT 0.072 0.153 0.218 0.171 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.5 0.243 ;

	END

END NOR2x2_ASAP7_75t_R

MACRO NOR2xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR2xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.143 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.094 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NOR2xp33_ASAP7_75t_R

MACRO NOR2xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR2xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.127 0.095 0.145 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.063 0.163 0.081 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END NOR2xp67_ASAP7_75t_R

MACRO NOR3x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR3x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.202 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.153 0.468 0.171 ;
			RECT 0.45 0.063 0.468 0.171 ;
			RECT 0.396 0.063 0.468 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.153 0.306 0.171 ;
			RECT 0.288 0.063 0.306 0.171 ;
			RECT 0.234 0.063 0.306 0.081 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.225 0.5 0.243 ;
			RECT 0.094 0.189 0.338 0.207 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END NOR3x1_ASAP7_75t_R

MACRO NOR3x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR3x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.904 0.189 1.062 0.207 ;
			RECT 1.044 0.027 1.062 0.207 ;
			RECT 0.018 0.027 1.062 0.045 ;
			RECT 0.018 0.189 0.176 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.169 0.072 0.908 0.09 ;
			LAYER M1 ;
			RECT 0.885 0.063 0.903 0.162 ;
			RECT 0.866 0.063 0.903 0.081 ;
			RECT 0.174 0.063 0.211 0.081 ;
			RECT 0.174 0.063 0.192 0.164 ;
			LAYER V1 ;
			RECT 0.174 0.072 0.192 0.09 ;
			RECT 0.885 0.072 0.903 0.09 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.725 0.063 0.743 0.164 ;
			RECT 0.338 0.063 0.743 0.081 ;
			RECT 0.338 0.063 0.356 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.547 0.106 0.565 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.742 0.225 0.986 0.243 ;
			RECT 0.256 0.189 0.824 0.207 ;
			RECT 0.418 0.225 0.662 0.243 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END NOR3x2_ASAP7_75t_R

MACRO NOR3xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR3xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.176 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END NOR3xp33_ASAP7_75t_R

MACRO NOR4xp25_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR4xp25_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.04 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END NOR4xp25_ASAP7_75t_R

MACRO NOR4xp75_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR4xp75_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.58 0.189 0.738 0.207 ;
			RECT 0.72 0.027 0.738 0.207 ;
			RECT 0.094 0.027 0.738 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.07 0.63 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.531 0.151 0.549 0.2 ;
			RECT 0.504 0.151 0.549 0.169 ;
			RECT 0.504 0.07 0.522 0.169 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.151 0.306 0.169 ;
			RECT 0.288 0.07 0.306 0.169 ;
			RECT 0.207 0.151 0.225 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.057 0.243 ;
			RECT 0.018 0.027 0.057 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.412 0.225 0.666 0.243 ;
			RECT 0.256 0.189 0.499 0.207 ;
			RECT 0.092 0.225 0.34 0.243 ;

	END

END NOR4xp75_ASAP7_75t_R

MACRO NOR5xp2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN NOR5xp2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.017 0.027 0.338 0.045 ;
			RECT 0.017 0.225 0.07 0.243 ;
			RECT 0.017 0.027 0.037 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END NOR5xp2_ASAP7_75t_R

MACRO O2A1O1Ixp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN O2A1O1Ixp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.206 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.225 0.243 ;
			RECT 0.04 0.063 0.176 0.081 ;

	END

END O2A1O1Ixp33_ASAP7_75t_R

MACRO O2A1O1Ixp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN O2A1O1Ixp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.315 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.252 0.164 ;
			RECT 0.072 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.189 0.338 0.207 ;
			RECT 0.148 0.027 0.279 0.045 ;
			RECT 0.094 0.225 0.23 0.243 ;

	END

END O2A1O1Ixp5_ASAP7_75t_R

MACRO OA211x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA211x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.296 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.286 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.234 0.189 0.306 0.207 ;
			RECT 0.288 0.063 0.306 0.207 ;
			RECT 0.099 0.063 0.306 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OA211x2_ASAP7_75t_R

MACRO OA21x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA21x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.256 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.153 0.239 0.171 ;
			RECT 0.18 0.106 0.198 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.225 0.224 0.243 ;
			RECT 0.206 0.189 0.224 0.243 ;
			RECT 0.206 0.189 0.306 0.207 ;
			RECT 0.288 0.063 0.306 0.207 ;
			RECT 0.099 0.063 0.306 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OA21x2_ASAP7_75t_R

MACRO OA221x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA221x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.225 0.117 0.243 ;
			RECT 0.099 0.189 0.117 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.099 0.252 0.207 ;
			RECT 0.215 0.099 0.252 0.117 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.593 0.189 0.63 0.207 ;
			RECT 0.612 0.099 0.63 0.207 ;
			RECT 0.593 0.099 0.63 0.117 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.099 0.522 0.207 ;
			RECT 0.485 0.099 0.522 0.117 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.72 0.189 0.757 0.207 ;
			RECT 0.72 0.099 0.757 0.117 ;
			RECT 0.72 0.099 0.738 0.207 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.144 0.225 0.846 0.243 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.144 0.126 0.162 0.243 ;
			RECT 0.121 0.126 0.162 0.144 ;
			RECT 0.741 0.063 0.846 0.081 ;
			RECT 0.472 0.027 0.824 0.045 ;
			RECT 0.202 0.063 0.668 0.081 ;

	END

END OA221x2_ASAP7_75t_R

MACRO OA222x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA222x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.531 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.526 0.027 0.63 0.045 ;
			RECT 0.531 0.189 0.549 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.009 0.225 0.504 0.243 ;
			RECT 0.486 0.126 0.504 0.243 ;
			RECT 0.009 0.063 0.027 0.243 ;
			RECT 0.486 0.126 0.554 0.144 ;
			RECT 0.009 0.063 0.122 0.081 ;
			RECT 0.202 0.063 0.36 0.081 ;
			RECT 0.342 0.027 0.36 0.081 ;
			RECT 0.342 0.027 0.468 0.045 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OA222x2_ASAP7_75t_R

MACRO OA22x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA22x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.071 0.225 0.122 0.243 ;
			RECT 0.071 0.027 0.122 0.045 ;
			RECT 0.071 0.027 0.091 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.236 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.063 0.414 0.2 ;
			RECT 0.367 0.063 0.414 0.081 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.18 0.225 0.392 0.243 ;
			RECT 0.18 0.063 0.198 0.243 ;
			RECT 0.137 0.126 0.198 0.144 ;
			RECT 0.18 0.063 0.333 0.081 ;
			RECT 0.256 0.027 0.5 0.045 ;

	END

END OA22x2_ASAP7_75t_R

MACRO OA31x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA31x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.693 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.053 0.189 0.09 0.207 ;
			RECT 0.072 0.099 0.09 0.207 ;
			RECT 0.053 0.099 0.09 0.117 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.126 0.189 0.163 0.207 ;
			RECT 0.126 0.106 0.144 0.207 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.126 0.414 0.144 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.323 0.063 0.36 0.081 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.153 0.522 0.171 ;
			RECT 0.504 0.106 0.522 0.171 ;

		END 

	END B1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.369 0.189 0.576 0.207 ;
			RECT 0.558 0.063 0.576 0.207 ;
			RECT 0.558 0.126 0.667 0.144 ;
			RECT 0.418 0.063 0.576 0.081 ;
			RECT 0.317 0.225 0.446 0.243 ;
			RECT 0.317 0.189 0.335 0.243 ;
			RECT 0.202 0.189 0.335 0.207 ;
			RECT 0.094 0.027 0.5 0.045 ;
			RECT 0.04 0.063 0.284 0.081 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END OA31x2_ASAP7_75t_R

MACRO OA331x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA331x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.166 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.099 0.186 0.117 0.243 ;
			RECT 0.072 0.186 0.117 0.204 ;
			RECT 0.072 0.115 0.09 0.204 ;
			RECT 0.471 0.063 0.522 0.081 ;
			RECT 0.234 0.063 0.393 0.081 ;
			RECT 0.234 0.027 0.252 0.081 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.308 0.027 0.447 0.045 ;

	END

END OA331x1_ASAP7_75t_R

MACRO OA331x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA331x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.045 0.225 0.122 0.243 ;
			RECT 0.045 0.027 0.122 0.045 ;
			RECT 0.045 0.027 0.063 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.166 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.153 0.186 0.171 0.243 ;
			RECT 0.126 0.186 0.171 0.204 ;
			RECT 0.126 0.115 0.144 0.204 ;
			RECT 0.525 0.063 0.576 0.081 ;
			RECT 0.288 0.063 0.447 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.202 0.027 0.306 0.045 ;
			RECT 0.362 0.027 0.501 0.045 ;

	END

END OA331x2_ASAP7_75t_R

MACRO OA332x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA332x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.094 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.126 0.189 0.144 0.243 ;
			RECT 0.072 0.189 0.144 0.207 ;
			RECT 0.072 0.119 0.09 0.207 ;
			RECT 0.471 0.063 0.576 0.081 ;
			RECT 0.234 0.063 0.393 0.081 ;
			RECT 0.234 0.027 0.252 0.081 ;
			RECT 0.146 0.027 0.252 0.045 ;
			RECT 0.308 0.027 0.556 0.045 ;

	END

END OA332x1_ASAP7_75t_R

MACRO OA332x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA332x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.137 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.18 0.225 0.63 0.243 ;
			RECT 0.612 0.063 0.63 0.243 ;
			RECT 0.18 0.189 0.198 0.243 ;
			RECT 0.126 0.189 0.198 0.207 ;
			RECT 0.126 0.119 0.144 0.207 ;
			RECT 0.525 0.063 0.63 0.081 ;
			RECT 0.288 0.063 0.447 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.2 0.027 0.306 0.045 ;
			RECT 0.362 0.027 0.61 0.045 ;

	END

END OA332x2_ASAP7_75t_R

MACRO OA333x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA333x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.63 0.243 ;
			RECT 0.612 0.063 0.63 0.243 ;
			RECT 0.099 0.186 0.117 0.243 ;
			RECT 0.072 0.186 0.117 0.204 ;
			RECT 0.072 0.115 0.09 0.204 ;
			RECT 0.467 0.063 0.63 0.081 ;
			RECT 0.232 0.063 0.394 0.081 ;
			RECT 0.232 0.027 0.25 0.081 ;
			RECT 0.147 0.027 0.25 0.045 ;
			RECT 0.309 0.027 0.569 0.045 ;

	END

END OA333x1_ASAP7_75t_R

MACRO OA333x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA333x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 0.122 0.243 ;
			RECT 0.072 0.027 0.122 0.045 ;
			RECT 0.072 0.027 0.09 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.106 0.63 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.684 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.153 0.186 0.171 0.243 ;
			RECT 0.126 0.186 0.171 0.204 ;
			RECT 0.126 0.115 0.144 0.204 ;
			RECT 0.521 0.063 0.684 0.081 ;
			RECT 0.286 0.063 0.448 0.081 ;
			RECT 0.286 0.027 0.304 0.081 ;
			RECT 0.201 0.027 0.304 0.045 ;
			RECT 0.363 0.027 0.623 0.045 ;

	END

END OA333x2_ASAP7_75t_R

MACRO OA33x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OA33x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.225 0.117 0.243 ;
			RECT 0.099 0.189 0.117 0.243 ;
			RECT 0.062 0.189 0.117 0.207 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.144 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.144 0.126 0.162 0.243 ;
			RECT 0.121 0.126 0.162 0.144 ;
			RECT 0.364 0.063 0.522 0.081 ;
			RECT 0.202 0.027 0.446 0.045 ;

	END

END OA33x2_ASAP7_75t_R

MACRO OAI211xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI211xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.099 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI211xp5_ASAP7_75t_R

MACRO OAI21x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI21x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.369 0.027 0.414 0.045 ;
			RECT 0.018 0.027 0.063 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.189 0.306 0.207 ;
			RECT 0.288 0.106 0.306 0.207 ;
			RECT 0.126 0.106 0.144 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.19 0.127 0.256 0.145 ;
			RECT 0.19 0.099 0.227 0.171 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.072 0.063 0.36 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.027 0.333 0.045 ;

	END

END OAI21x1_ASAP7_75t_R

MACRO OAI21xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI21xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.099 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.203 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI21xp33_ASAP7_75t_R

MACRO OAI21xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI21xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.099 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.203 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI21xp5_ASAP7_75t_R

MACRO OAI221xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI221xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.23 0.243 ;
			RECT 0.018 0.063 0.123 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.201 0.063 0.339 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI221xp5_ASAP7_75t_R

MACRO OAI222xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI222xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.522 0.243 ;
			RECT 0.504 0.055 0.522 0.243 ;
			RECT 0.018 0.063 0.122 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.063 0.36 0.081 ;
			RECT 0.342 0.027 0.36 0.081 ;
			RECT 0.342 0.027 0.468 0.045 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI222xp33_ASAP7_75t_R

MACRO OAI22x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI22x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.038 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.309 0.063 0.522 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.153 0.379 0.171 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.189 0.468 0.207 ;
			RECT 0.45 0.099 0.468 0.207 ;
			RECT 0.431 0.099 0.468 0.117 ;
			RECT 0.288 0.118 0.306 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.161 0.153 0.198 0.171 ;
			RECT 0.18 0.063 0.198 0.171 ;
			RECT 0.161 0.063 0.198 0.081 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.189 0.252 0.207 ;
			RECT 0.234 0.116 0.252 0.207 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.207 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.5 0.045 ;

	END

END OAI22x1_ASAP7_75t_R

MACRO OAI22xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI22xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.063 0.117 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.225 0.275 0.243 ;
			RECT 0.234 0.07 0.252 0.243 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI22xp33_ASAP7_75t_R

MACRO OAI22xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI22xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.063 0.117 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.225 0.275 0.243 ;
			RECT 0.234 0.07 0.252 0.243 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.063 0.198 0.164 ;
			RECT 0.151 0.063 0.198 0.081 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI22xp5_ASAP7_75t_R

MACRO OAI311xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI311xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.198 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END B1
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.027 0.234 0.045 ;

	END

END OAI311xp33_ASAP7_75t_R

MACRO OAI31xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI31xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.256 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.093 0.027 0.23 0.045 ;

	END

END OAI31xp33_ASAP7_75t_R

MACRO OAI31xp67_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI31xp67_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.063 0.663 0.081 ;
			RECT 0.202 0.189 0.252 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.666 0.126 0.684 0.198 ;
			RECT 0.553 0.126 0.684 0.144 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.126 0.419 0.144 ;
			RECT 0.288 0.126 0.306 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.225 0.663 0.243 ;
			RECT 0.364 0.189 0.608 0.207 ;
			RECT 0.04 0.027 0.554 0.045 ;
			RECT 0.094 0.225 0.446 0.243 ;

	END

END OAI31xp67_ASAP7_75t_R

MACRO OAI321xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI321xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.198 0.225 0.414 0.243 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.31 0.063 0.414 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.396 0.045 ;
			RECT 0.094 0.063 0.23 0.081 ;

	END

END OAI321xp33_ASAP7_75t_R

MACRO OAI322xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI322xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.147 0.225 0.468 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.364 0.063 0.468 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.105 0.306 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.105 0.36 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.027 0.45 0.045 ;
			RECT 0.039 0.063 0.284 0.081 ;

	END

END OAI322xp33_ASAP7_75t_R

MACRO OAI32xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI32xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.36 0.243 ;
			RECT 0.342 0.063 0.36 0.243 ;
			RECT 0.256 0.063 0.36 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.063 0.222 0.081 ;
			RECT 0.18 0.063 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.027 0.338 0.045 ;

	END

END OAI32xp33_ASAP7_75t_R

MACRO OAI331xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI331xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.468 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.417 0.063 0.468 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.393 0.045 ;
			RECT 0.092 0.063 0.339 0.081 ;

	END

END OAI331xp33_ASAP7_75t_R

MACRO OAI332xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI332xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.417 0.063 0.522 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.502 0.045 ;
			RECT 0.092 0.063 0.339 0.081 ;

	END

END OAI332xp33_ASAP7_75t_R

MACRO OAI333xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI333xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.413 0.063 0.576 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.515 0.045 ;
			RECT 0.094 0.063 0.34 0.081 ;

	END

END OAI333xp33_ASAP7_75t_R

MACRO OAI33xp33_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OAI33xp33_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.414 0.243 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.256 0.063 0.414 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.092 0.027 0.338 0.045 ;

	END

END OAI33xp33_ASAP7_75t_R

MACRO OR2x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR2x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.207 0.027 0.306 0.045 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.077 0.144 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.186 0.243 ;
			RECT 0.168 0.027 0.186 0.243 ;
			RECT 0.168 0.126 0.227 0.144 ;
			RECT 0.094 0.027 0.186 0.045 ;

	END

END OR2x2_ASAP7_75t_R

MACRO OR2x4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR2x4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.207 0.027 0.414 0.045 ;
			RECT 0.315 0.184 0.333 0.243 ;
			RECT 0.315 0.027 0.333 0.086 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.077 0.144 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.187 0.243 ;
			RECT 0.169 0.027 0.187 0.243 ;
			RECT 0.169 0.126 0.227 0.144 ;
			RECT 0.094 0.027 0.187 0.045 ;

	END

END OR2x4_ASAP7_75t_R

MACRO OR2x6_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR2x6_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.31 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.063 0.144 0.122 ;
			RECT 0.018 0.063 0.144 0.081 ;
			RECT 0.018 0.063 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.153 0.252 0.171 ;
			RECT 0.234 0.121 0.252 0.171 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.189 0.306 0.207 ;
			RECT 0.288 0.07 0.306 0.207 ;
			RECT 0.234 0.07 0.306 0.088 ;
			RECT 0.234 0.027 0.252 0.088 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END OR2x6_ASAP7_75t_R

MACRO OR3x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR3x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.183 0.306 0.201 ;
			RECT 0.288 0.076 0.306 0.201 ;
			RECT 0.261 0.076 0.306 0.094 ;
			RECT 0.261 0.183 0.279 0.235 ;
			RECT 0.261 0.034 0.279 0.094 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.262 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END OR3x1_ASAP7_75t_R

MACRO OR3x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR3x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.261 0.027 0.36 0.045 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.24 0.243 ;
			RECT 0.222 0.027 0.24 0.243 ;
			RECT 0.222 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.24 0.045 ;

	END

END OR3x2_ASAP7_75t_R

MACRO OR3x4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR3x4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.261 0.027 0.468 0.045 ;
			RECT 0.369 0.184 0.387 0.243 ;
			RECT 0.369 0.027 0.387 0.086 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.241 0.243 ;
			RECT 0.223 0.027 0.241 0.243 ;
			RECT 0.223 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.241 0.045 ;

	END

END OR3x4_ASAP7_75t_R

MACRO OR4x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR4x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.072 0.066 0.09 0.152 ;
			RECT 0.072 0.066 0.117 0.084 ;
			RECT 0.099 0.027 0.117 0.084 ;
			RECT 0.099 0.027 0.36 0.045 ;

	END

END OR4x1_ASAP7_75t_R

MACRO OR4x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR4x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.364 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.099 0.063 0.117 0.149 ;
			RECT 0.099 0.063 0.171 0.081 ;
			RECT 0.153 0.027 0.171 0.081 ;
			RECT 0.153 0.027 0.414 0.045 ;

	END

END OR4x2_ASAP7_75t_R

MACRO OR5x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR5x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.35 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.349 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.07 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.288 0.063 0.36 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.018 0.027 0.306 0.045 ;

	END

END OR5x1_ASAP7_75t_R

MACRO OR5x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN OR5x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.343 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.07 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.288 0.063 0.36 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.018 0.027 0.306 0.045 ;

	END

END OR5x2_ASAP7_75t_R

MACRO SDFHx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFHx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.332 0.243 ;
			RECT 1.314 0.027 1.332 0.243 ;
			RECT 1.282 0.027 1.332 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.185 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.185 0.117 0.203 ;
			RECT 0.072 0.081 0.09 0.203 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.284 0.108 0.436 0.126 ;
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.164 ;
			LAYER V1 ;
			RECT 0.396 0.108 0.414 0.126 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.467 0.108 0.59 0.126 ;
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;
			LAYER V1 ;
			RECT 0.504 0.108 0.522 0.126 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.797 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.021 0.225 0.068 0.243 ;
			RECT 0.021 0.027 0.039 0.243 ;
			RECT 0.021 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.016 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.021 0.144 0.039 0.162 ;

	END

END SDFHx1_ASAP7_75t_R

MACRO SDFHx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFHx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.282 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.019 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx2_ASAP7_75t_R

MACRO SDFHx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFHx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.458 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.44 0.243 ;
			RECT 1.422 0.027 1.44 0.243 ;
			RECT 1.282 0.027 1.44 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.458 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.458 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.019 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx3_ASAP7_75t_R

MACRO SDFHx4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFHx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.674 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.444 0.225 1.656 0.243 ;
			RECT 1.637 0.027 1.656 0.243 ;
			RECT 1.444 0.027 1.656 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.164 ;
			RECT 0.378 0.225 0.459 0.243 ;
			RECT 0.378 0.099 0.468 0.117 ;
			RECT 0.378 0.099 0.396 0.243 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.599 0.081 ;
			RECT 0.558 0.063 0.576 0.164 ;
			RECT 0.234 0.126 0.289 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;
			LAYER V1 ;
			RECT 0.234 0.072 0.252 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.027 0.767 0.045 ;
			RECT 0.639 0.063 0.711 0.081 ;
			RECT 0.693 0.027 0.711 0.081 ;
			RECT 0.612 0.106 0.657 0.124 ;
			RECT 0.639 0.063 0.657 0.124 ;
			RECT 0.612 0.106 0.63 0.164 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.674 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.674 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.059 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.368 0.126 1.447 0.144 ;
			RECT 1.242 0.126 1.283 0.144 ;
			RECT 1.242 0.027 1.26 0.144 ;
			RECT 1.113 0.027 1.386 0.045 ;
			RECT 1.206 0.182 1.332 0.2 ;
			RECT 1.314 0.081 1.332 0.2 ;
			RECT 1.206 0.106 1.224 0.2 ;
			RECT 1.287 0.081 1.332 0.099 ;
			RECT 0.882 0.063 0.9 0.164 ;
			RECT 0.882 0.063 0.981 0.081 ;
			RECT 0.801 0.225 0.954 0.243 ;
			RECT 0.936 0.106 0.954 0.243 ;
			RECT 0.801 0.189 0.819 0.243 ;
			RECT 0.738 0.189 0.819 0.207 ;
			RECT 0.738 0.07 0.756 0.207 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.504 0.063 0.522 0.164 ;
			RECT 0.342 0.063 0.522 0.081 ;
			RECT 0.31 0.027 0.36 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.126 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.09 0.045 ;
			RECT 1.152 0.106 1.17 0.2 ;
			RECT 1.098 0.07 1.116 0.164 ;
			RECT 1.044 0.106 1.062 0.2 ;
			RECT 0.828 0.07 0.846 0.167 ;
			RECT 0.774 0.07 0.792 0.164 ;
			RECT 0.58 0.225 0.77 0.243 ;
			RECT 0.684 0.121 0.702 0.167 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.423 0.189 0.662 0.207 ;
			RECT 0.126 0.106 0.144 0.2 ;
			LAYER M2 ;
			RECT 0.019 0.144 1.175 0.162 ;
			RECT 0.175 0.108 1.121 0.126 ;
			LAYER V1 ;
			RECT 1.152 0.144 1.17 0.162 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 1.044 0.144 1.062 0.162 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.108 0.792 0.126 ;
			RECT 0.684 0.144 0.702 0.162 ;
			RECT 0.18 0.108 0.198 0.126 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx4_ASAP7_75t_R

MACRO SDFLx1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFLx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.332 0.243 ;
			RECT 1.314 0.027 1.332 0.243 ;
			RECT 1.282 0.027 1.332 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.797 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx1_ASAP7_75t_R

MACRO SDFLx2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFLx2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.282 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx2_ASAP7_75t_R

MACRO SDFLx3_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFLx3_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.458 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.44 0.243 ;
			RECT 1.422 0.027 1.44 0.243 ;
			RECT 1.282 0.027 1.44 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.458 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.458 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx3_ASAP7_75t_R

MACRO SDFLx4_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN SDFLx4_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.674 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.444 0.225 1.656 0.243 ;
			RECT 1.637 0.027 1.656 0.243 ;
			RECT 1.444 0.027 1.656 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.164 ;
			RECT 0.378 0.225 0.459 0.243 ;
			RECT 0.378 0.099 0.468 0.117 ;
			RECT 0.378 0.099 0.396 0.243 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.599 0.081 ;
			RECT 0.558 0.063 0.576 0.164 ;
			RECT 0.234 0.126 0.289 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;
			LAYER V1 ;
			RECT 0.234 0.072 0.252 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.027 0.767 0.045 ;
			RECT 0.639 0.063 0.711 0.081 ;
			RECT 0.693 0.027 0.711 0.081 ;
			RECT 0.612 0.106 0.657 0.124 ;
			RECT 0.639 0.063 0.657 0.124 ;
			RECT 0.612 0.106 0.63 0.164 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.674 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.674 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.059 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.368 0.126 1.447 0.144 ;
			RECT 1.242 0.126 1.283 0.144 ;
			RECT 1.242 0.027 1.26 0.144 ;
			RECT 1.113 0.027 1.386 0.045 ;
			RECT 1.206 0.182 1.332 0.2 ;
			RECT 1.314 0.081 1.332 0.2 ;
			RECT 1.206 0.106 1.224 0.2 ;
			RECT 1.287 0.081 1.332 0.099 ;
			RECT 0.882 0.063 0.9 0.164 ;
			RECT 0.882 0.063 0.981 0.081 ;
			RECT 0.801 0.225 0.954 0.243 ;
			RECT 0.936 0.106 0.954 0.243 ;
			RECT 0.801 0.189 0.819 0.243 ;
			RECT 0.738 0.189 0.819 0.207 ;
			RECT 0.738 0.07 0.756 0.207 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.504 0.063 0.522 0.164 ;
			RECT 0.342 0.063 0.522 0.081 ;
			RECT 0.31 0.027 0.36 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.126 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.108 0.047 0.126 ;
			RECT 0.009 0.027 0.09 0.045 ;
			RECT 1.152 0.106 1.17 0.2 ;
			RECT 1.098 0.07 1.116 0.164 ;
			RECT 1.044 0.106 1.062 0.2 ;
			RECT 0.828 0.07 0.846 0.167 ;
			RECT 0.774 0.07 0.792 0.164 ;
			RECT 0.58 0.225 0.77 0.243 ;
			RECT 0.684 0.121 0.702 0.167 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.423 0.189 0.662 0.207 ;
			RECT 0.126 0.103 0.144 0.2 ;
			LAYER M2 ;
			RECT 0.175 0.144 1.175 0.162 ;
			RECT 0.019 0.108 1.121 0.126 ;
			LAYER V1 ;
			RECT 1.152 0.144 1.17 0.162 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 1.044 0.144 1.062 0.162 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.108 0.792 0.126 ;
			RECT 0.684 0.144 0.702 0.162 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.108 0.144 0.126 ;
			RECT 0.024 0.108 0.042 0.126 ;

	END

END SDFLx4_ASAP7_75t_R

MACRO TAPCELL_ASAP7_75t_R
	CLASS CORE WELLTAP ;
	FOREIGN TAPCELL_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.108 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.108 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.108 0.279 ;

		END 

	END VDD

END TAPCELL_ASAP7_75t_R

MACRO TAPCELL_WITH_FILLER_ASAP7_75t_R
	CLASS CORE WELLTAP ;
	FOREIGN TAPCELL_WITH_FILLER_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END TAPCELL_WITH_FILLER_ASAP7_75t_R

MACRO TIEHIx1_ASAP7_75t_R
	CLASS CORE TIEHIGH ;
	FOREIGN TIEHIx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN H
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.07 0.144 0.243 ;
			RECT 0.067 0.07 0.144 0.088 ;

		END 

	END H
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.155 0.095 0.173 ;
			RECT 0.018 0.027 0.036 0.173 ;
			RECT 0.018 0.027 0.068 0.045 ;

	END

END TIEHIx1_ASAP7_75t_R

MACRO TIELOx1_ASAP7_75t_R
	CLASS CORE TIELOW ;
	FOREIGN TIELOx1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN L
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.067 0.182 0.144 0.2 ;
			RECT 0.126 0.027 0.144 0.2 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END L
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.097 0.036 0.243 ;
			RECT 0.018 0.097 0.095 0.115 ;

	END

END TIELOx1_ASAP7_75t_R

MACRO XNOR2x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN XNOR2x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.612 0.243 ;
			RECT 0.45 0.077 0.468 0.243 ;
			RECT 0.418 0.077 0.468 0.095 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.121 0.18 0.581 0.198 ;
			LAYER M1 ;
			RECT 0.526 0.189 0.576 0.207 ;
			RECT 0.558 0.121 0.576 0.207 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			LAYER V1 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.558 0.18 0.576 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.298 0.072 0.527 0.09 ;
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.152 ;
			RECT 0.305 0.126 0.365 0.144 ;
			RECT 0.305 0.067 0.323 0.144 ;
			RECT 0.213 0.067 0.323 0.085 ;
			RECT 0.213 0.027 0.231 0.085 ;
			RECT 0.018 0.027 0.231 0.045 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.027 0.036 0.236 ;
			LAYER V1 ;
			RECT 0.305 0.072 0.323 0.09 ;
			RECT 0.504 0.072 0.522 0.09 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.092 0.225 0.193 0.243 ;
			RECT 0.174 0.189 0.193 0.243 ;
			RECT 0.174 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.174 0.082 0.192 0.243 ;
			RECT 0.256 0.027 0.608 0.045 ;

	END

END XNOR2x1_ASAP7_75t_R

MACRO XNOR2x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN XNOR2x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.472 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.44 0.243 ;
			RECT 0.422 0.126 0.44 0.243 ;
			RECT 0.391 0.126 0.44 0.144 ;
			RECT 0.261 0.183 0.279 0.243 ;
			RECT 0.126 0.183 0.279 0.201 ;
			RECT 0.126 0.12 0.144 0.201 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.189 0.38 0.207 ;
			RECT 0.342 0.107 0.36 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.063 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.477 0.063 0.495 0.151 ;
			RECT 0.423 0.063 0.495 0.081 ;
			RECT 0.423 0.027 0.441 0.081 ;
			RECT 0.018 0.027 0.441 0.045 ;
			RECT 0.302 0.063 0.32 0.195 ;
			RECT 0.072 0.063 0.09 0.149 ;
			RECT 0.072 0.063 0.392 0.081 ;
			RECT 0.099 0.225 0.23 0.243 ;

	END

END XNOR2x2_ASAP7_75t_R

MACRO XNOR2xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN XNOR2xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.423 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.207 0.063 0.36 0.081 ;
			RECT 0.207 0.027 0.225 0.081 ;
			RECT 0.072 0.027 0.225 0.045 ;
			RECT 0.072 0.027 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.075 0.18 0.243 ;
			RECT 0.162 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.261 0.027 0.387 0.045 ;

	END

END XNOR2xp5_ASAP7_75t_R

MACRO XOR2x1_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN XOR2x1_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.027 0.612 0.045 ;
			RECT 0.418 0.175 0.468 0.193 ;
			RECT 0.45 0.027 0.468 0.193 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.298 0.18 0.527 0.198 ;
			LAYER M1 ;
			RECT 0.504 0.118 0.522 0.2 ;
			RECT 0.305 0.126 0.365 0.144 ;
			RECT 0.213 0.185 0.323 0.203 ;
			RECT 0.305 0.126 0.323 0.203 ;
			RECT 0.018 0.225 0.231 0.243 ;
			RECT 0.213 0.185 0.231 0.243 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.243 ;
			LAYER V1 ;
			RECT 0.305 0.18 0.323 0.198 ;
			RECT 0.504 0.18 0.522 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.121 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.576 0.149 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.126 0.063 0.144 0.149 ;
			RECT 0.107 0.063 0.144 0.081 ;
			LAYER V1 ;
			RECT 0.126 0.072 0.144 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.174 0.027 0.192 0.188 ;
			RECT 0.396 0.063 0.414 0.149 ;
			RECT 0.174 0.063 0.414 0.081 ;
			RECT 0.174 0.027 0.193 0.081 ;
			RECT 0.092 0.027 0.193 0.045 ;
			RECT 0.256 0.225 0.608 0.243 ;

	END

END XOR2x1_ASAP7_75t_R

MACRO XOR2x2_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN XOR2x2_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.472 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.38 0.081 ;
			RECT 0.342 0.063 0.36 0.163 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.422 0.027 0.44 0.163 ;
			RECT 0.391 0.126 0.44 0.144 ;
			RECT 0.261 0.027 0.44 0.045 ;
			RECT 0.126 0.069 0.279 0.087 ;
			RECT 0.261 0.027 0.279 0.087 ;
			RECT 0.126 0.069 0.144 0.15 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.441 0.243 ;
			RECT 0.423 0.189 0.441 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.423 0.189 0.495 0.207 ;
			RECT 0.477 0.119 0.495 0.207 ;
			RECT 0.018 0.027 0.063 0.045 ;
			RECT 0.072 0.189 0.392 0.207 ;
			RECT 0.302 0.075 0.32 0.207 ;
			RECT 0.072 0.121 0.09 0.207 ;
			RECT 0.099 0.027 0.23 0.045 ;

	END

END XOR2x2_ASAP7_75t_R

MACRO XOR2xp5_ASAP7_75t_R
	CLASS CORE ;
	FOREIGN XOR2xp5_ASAP7_75t_R 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.423 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.256 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.189 0.36 0.207 ;
			RECT 0.342 0.12 0.36 0.207 ;
			RECT 0.018 0.225 0.225 0.243 ;
			RECT 0.207 0.189 0.225 0.243 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.106 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.162 0.027 0.18 0.195 ;
			RECT 0.396 0.063 0.414 0.149 ;
			RECT 0.162 0.063 0.414 0.081 ;
			RECT 0.094 0.027 0.18 0.045 ;
			RECT 0.256 0.225 0.387 0.243 ;

	END

END XOR2xp5_ASAP7_75t_R

MACRO A2O1A1Ixp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN A2O1A1Ixp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.214 0.215 0.306 0.233 ;
			RECT 0.288 0.037 0.306 0.233 ;
			RECT 0.262 0.037 0.306 0.055 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.081 0.252 0.19 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.23 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END A2O1A1Ixp33_ASAP7_75t_L

MACRO A2O1A1O1Ixp25_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN A2O1A1O1Ixp25_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.423 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.261 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.127 0.414 0.145 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.207 0.225 0.387 0.243 ;
			RECT 0.04 0.027 0.225 0.045 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END A2O1A1O1Ixp25_ASAP7_75t_L

MACRO AND2x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND2x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.207 0.027 0.306 0.045 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.027 0.18 0.243 ;
			RECT 0.162 0.126 0.203 0.144 ;
			RECT 0.07 0.027 0.088 0.086 ;
			RECT 0.07 0.027 0.18 0.045 ;

	END

END AND2x2_ASAP7_75t_L

MACRO AND2x4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND2x4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.31 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.028 0.252 0.15 ;
			RECT 0.072 0.028 0.252 0.046 ;
			RECT 0.072 0.028 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.107 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.231 0.243 ;
			RECT 0.18 0.064 0.198 0.243 ;
			RECT 0.179 0.182 0.306 0.2 ;
			RECT 0.288 0.121 0.306 0.2 ;
			RECT 0.115 0.064 0.198 0.082 ;

	END

END AND2x4_ASAP7_75t_L

MACRO AND2x6_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND2x6_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.554 0.243 ;
			RECT 0.31 0.027 0.554 0.045 ;
			RECT 0.45 0.027 0.468 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.028 0.252 0.15 ;
			RECT 0.072 0.028 0.252 0.046 ;
			RECT 0.072 0.028 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.107 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.231 0.243 ;
			RECT 0.18 0.064 0.198 0.243 ;
			RECT 0.179 0.182 0.306 0.2 ;
			RECT 0.288 0.121 0.306 0.2 ;
			RECT 0.115 0.064 0.198 0.082 ;

	END

END AND2x6_ASAP7_75t_L

MACRO AND3x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND3x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.183 0.306 0.201 ;
			RECT 0.288 0.076 0.306 0.201 ;
			RECT 0.261 0.076 0.306 0.094 ;
			RECT 0.261 0.183 0.279 0.235 ;
			RECT 0.261 0.034 0.279 0.094 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.263 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END AND3x1_ASAP7_75t_L

MACRO AND3x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND3x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.261 0.027 0.36 0.045 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END AND3x2_ASAP7_75t_L

MACRO AND3x4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND3x4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.23 0.243 ;
			RECT 0.018 0.027 0.23 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.189 0.649 0.207 ;
			RECT 0.612 0.099 0.649 0.117 ;
			RECT 0.612 0.099 0.63 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.189 0.541 0.207 ;
			RECT 0.504 0.099 0.541 0.117 ;
			RECT 0.504 0.099 0.522 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.26 0.225 0.746 0.243 ;
			RECT 0.728 0.027 0.746 0.243 ;
			RECT 0.26 0.042 0.278 0.243 ;
			RECT 0.218 0.126 0.278 0.144 ;
			RECT 0.634 0.027 0.746 0.045 ;
			RECT 0.472 0.063 0.701 0.081 ;
			RECT 0.31 0.027 0.554 0.045 ;

	END

END AND3x4_ASAP7_75t_L

MACRO AND4x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND4x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.299 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.164 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.234 0.189 0.306 0.207 ;
			RECT 0.288 0.12 0.306 0.207 ;
			RECT 0.018 0.027 0.085 0.045 ;

	END

END AND4x1_ASAP7_75t_L

MACRO AND4x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND4x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.164 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.153 0.189 0.171 0.243 ;
			RECT 0.099 0.189 0.171 0.207 ;
			RECT 0.099 0.119 0.117 0.207 ;
			RECT 0.364 0.027 0.414 0.045 ;

	END

END AND4x2_ASAP7_75t_L

MACRO AND5x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND5x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.349 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.35 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.164 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.288 0.189 0.36 0.207 ;
			RECT 0.342 0.116 0.36 0.207 ;
			RECT 0.018 0.027 0.07 0.045 ;

	END

END AND5x1_ASAP7_75t_L

MACRO AND5x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AND5x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.958 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.958 0.027 1.062 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.72 0.189 0.757 0.207 ;
			RECT 0.72 0.099 0.757 0.117 ;
			RECT 0.72 0.099 0.738 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.593 0.189 0.63 0.207 ;
			RECT 0.612 0.099 0.63 0.207 ;
			RECT 0.593 0.099 0.63 0.117 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.189 0.487 0.207 ;
			RECT 0.45 0.099 0.487 0.117 ;
			RECT 0.45 0.099 0.468 0.207 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.269 0.189 0.306 0.207 ;
			RECT 0.288 0.099 0.306 0.207 ;
			RECT 0.269 0.099 0.306 0.117 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.225 0.9 0.243 ;
			RECT 0.882 0.027 0.9 0.243 ;
			RECT 0.882 0.126 0.942 0.144 ;
			RECT 0.742 0.027 0.9 0.045 ;
			RECT 0.58 0.063 0.824 0.081 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.256 0.063 0.5 0.081 ;
			RECT 0.094 0.027 0.338 0.045 ;

	END

END AND5x2_ASAP7_75t_L

MACRO AO211x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO211x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.742 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.311 0.144 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.215 0.063 0.252 0.081 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.153 0.541 0.171 ;
			RECT 0.504 0.063 0.522 0.171 ;
			RECT 0.485 0.063 0.522 0.081 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.666 0.125 0.743 0.143 ;
			RECT 0.094 0.027 0.684 0.045 ;
			RECT 0.31 0.189 0.608 0.207 ;
			RECT 0.04 0.225 0.393 0.243 ;

	END

END AO211x2_ASAP7_75t_L

MACRO AO21x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO21x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.23 0.225 0.295 0.243 ;
			RECT 0.277 0.038 0.295 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.189 0.252 0.207 ;
			RECT 0.234 0.027 0.252 0.207 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AO21x1_ASAP7_75t_L

MACRO AO21x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO21x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.23 0.225 0.333 0.243 ;
			RECT 0.315 0.069 0.333 0.243 ;
			RECT 0.276 0.069 0.333 0.087 ;
			RECT 0.276 0.038 0.294 0.087 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.189 0.252 0.207 ;
			RECT 0.234 0.027 0.252 0.207 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AO21x2_ASAP7_75t_L

MACRO AO221x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO221x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.459 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.126 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;
			RECT 0.396 0.126 0.474 0.144 ;
			RECT 0.396 0.027 0.414 0.144 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.2 0.189 0.339 0.207 ;
			RECT 0.039 0.225 0.176 0.243 ;

	END

END AO221x1_ASAP7_75t_L

MACRO AO221x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO221x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.549 0.243 ;
			RECT 0.531 0.027 0.549 0.243 ;
			RECT 0.459 0.027 0.549 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.126 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;
			RECT 0.396 0.126 0.474 0.144 ;
			RECT 0.396 0.027 0.414 0.144 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.2 0.189 0.339 0.207 ;
			RECT 0.039 0.225 0.176 0.243 ;

	END

END AO221x2_ASAP7_75t_L

MACRO AO222x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO222x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.526 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.531 0.027 0.63 0.045 ;
			RECT 0.531 0.027 0.549 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.009 0.189 0.122 0.207 ;
			RECT 0.009 0.027 0.027 0.207 ;
			RECT 0.486 0.126 0.554 0.144 ;
			RECT 0.486 0.027 0.504 0.144 ;
			RECT 0.009 0.027 0.504 0.045 ;
			RECT 0.342 0.225 0.468 0.243 ;
			RECT 0.342 0.189 0.36 0.243 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO222x2_ASAP7_75t_L

MACRO AO22x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO22x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.418 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.287 0.081 ;
			RECT 0.234 0.063 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.342 0.126 0.419 0.144 ;
			RECT 0.107 0.027 0.36 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO22x1_ASAP7_75t_L

MACRO AO22x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO22x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.418 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.287 0.081 ;
			RECT 0.234 0.063 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.342 0.126 0.419 0.144 ;
			RECT 0.107 0.027 0.36 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO22x2_ASAP7_75t_L

MACRO AO31x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO31x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.741 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.742 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.099 0.576 0.149 ;
			RECT 0.504 0.099 0.576 0.117 ;
			RECT 0.485 0.153 0.522 0.171 ;
			RECT 0.504 0.099 0.522 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.414 0.149 ;
			RECT 0.288 0.099 0.414 0.117 ;
			RECT 0.288 0.153 0.325 0.171 ;
			RECT 0.288 0.07 0.306 0.171 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.059 0.207 ;
			RECT 0.018 0.027 0.059 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.612 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.612 0.189 0.63 0.243 ;
			RECT 0.199 0.189 0.63 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.666 0.126 0.797 0.144 ;
			RECT 0.2 0.063 0.252 0.081 ;
			RECT 0.526 0.027 0.684 0.045 ;
			RECT 0.364 0.063 0.608 0.081 ;
			RECT 0.04 0.225 0.554 0.243 ;
			RECT 0.094 0.027 0.447 0.045 ;

	END

END AO31x2_ASAP7_75t_L

MACRO AO322x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO322x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.634 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.634 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.153 0.325 0.171 ;
			RECT 0.288 0.063 0.325 0.081 ;
			RECT 0.288 0.063 0.306 0.171 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.063 0.541 0.081 ;
			RECT 0.504 0.063 0.522 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.396 0.189 0.576 0.207 ;
			RECT 0.558 0.126 0.576 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.558 0.126 0.743 0.144 ;
			RECT 0.04 0.027 0.446 0.045 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.189 0.198 0.243 ;
			RECT 0.18 0.189 0.338 0.207 ;
			RECT 0.256 0.225 0.5 0.243 ;

	END

END AO322x2_ASAP7_75t_L

MACRO AO32x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO32x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.063 0.063 0.081 ;
			RECT 0.045 0.034 0.063 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.062 0.126 0.108 0.144 ;
			RECT 0.09 0.027 0.108 0.144 ;
			RECT 0.09 0.027 0.414 0.045 ;
			RECT 0.148 0.225 0.392 0.243 ;

	END

END AO32x1_ASAP7_75t_L

MACRO AO32x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO32x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.068 0.117 0.086 ;
			RECT 0.099 0.037 0.117 0.086 ;
			RECT 0.018 0.068 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.189 0.33 0.207 ;
			RECT 0.288 0.07 0.306 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.364 0.189 0.468 0.207 ;
			RECT 0.45 0.027 0.468 0.207 ;
			RECT 0.093 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.468 0.045 ;
			RECT 0.202 0.225 0.446 0.243 ;

	END

END AO32x2_ASAP7_75t_L

MACRO AO331x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO331x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.081 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B3
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.072 0.063 0.09 0.152 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.522 0.045 ;
			RECT 0.308 0.189 0.447 0.207 ;
			RECT 0.146 0.225 0.393 0.243 ;

	END

END AO331x1_ASAP7_75t_L

MACRO AO331x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO331x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.027 0.135 0.045 ;
			RECT 0.072 0.225 0.122 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.126 0.063 0.144 0.152 ;
			RECT 0.126 0.063 0.198 0.081 ;
			RECT 0.18 0.027 0.198 0.081 ;
			RECT 0.18 0.027 0.576 0.045 ;
			RECT 0.362 0.189 0.501 0.207 ;
			RECT 0.2 0.225 0.447 0.243 ;

	END

END AO331x2_ASAP7_75t_L

MACRO AO332x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO332x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.094 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.072 0.063 0.09 0.151 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.576 0.045 ;
			RECT 0.146 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.234 0.189 0.393 0.207 ;
			RECT 0.308 0.225 0.556 0.243 ;

	END

END AO332x1_ASAP7_75t_L

MACRO AO332x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO332x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.148 0.045 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.189 0.63 0.207 ;
			RECT 0.612 0.027 0.63 0.207 ;
			RECT 0.126 0.063 0.144 0.151 ;
			RECT 0.126 0.063 0.198 0.081 ;
			RECT 0.18 0.027 0.198 0.081 ;
			RECT 0.18 0.027 0.63 0.045 ;
			RECT 0.2 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.288 0.189 0.447 0.207 ;
			RECT 0.362 0.225 0.61 0.243 ;

	END

END AO332x2_ASAP7_75t_L

MACRO AO333x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO333x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.081 0.045 ;
			RECT 0.018 0.225 0.069 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.063 0.09 0.152 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.63 0.045 ;
			RECT 0.31 0.189 0.576 0.207 ;
			RECT 0.148 0.225 0.395 0.243 ;

	END

END AO333x1_ASAP7_75t_L

MACRO AO333x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO333x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.081 0.117 0.099 ;
			RECT 0.099 0.045 0.117 0.099 ;
			RECT 0.018 0.081 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.07 0.63 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.067 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.684 0.045 ;
			RECT 0.364 0.189 0.63 0.207 ;
			RECT 0.202 0.225 0.449 0.243 ;

	END

END AO333x2_ASAP7_75t_L

MACRO AO33x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AO33x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.068 0.117 0.086 ;
			RECT 0.099 0.037 0.117 0.086 ;
			RECT 0.018 0.068 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.361 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.067 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.522 0.045 ;
			RECT 0.199 0.225 0.449 0.243 ;

	END

END AO33x2_ASAP7_75t_L

MACRO AOI211x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI211x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.519 0.189 0.63 0.207 ;
			RECT 0.612 0.027 0.63 0.207 ;
			RECT 0.091 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.126 0.229 0.144 ;
			RECT 0.18 0.189 0.223 0.207 ;
			RECT 0.18 0.063 0.22 0.081 ;
			RECT 0.18 0.063 0.198 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.123 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.153 0.442 0.171 ;
			RECT 0.396 0.063 0.442 0.081 ;
			RECT 0.396 0.063 0.414 0.171 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.126 0.554 0.144 ;
			RECT 0.504 0.063 0.55 0.081 ;
			RECT 0.504 0.063 0.522 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.288 0.189 0.449 0.207 ;
			RECT 0.361 0.225 0.608 0.243 ;

	END

END AOI211x1_ASAP7_75t_L

MACRO AOI211xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI211xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.04 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AOI211xp5_ASAP7_75t_L

MACRO AOI21x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI21x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.369 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.018 0.225 0.063 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.063 0.306 0.164 ;
			RECT 0.126 0.063 0.306 0.081 ;
			RECT 0.126 0.063 0.144 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.19 0.125 0.256 0.143 ;
			RECT 0.19 0.099 0.227 0.171 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.189 0.36 0.207 ;
			RECT 0.342 0.116 0.36 0.207 ;
			RECT 0.072 0.07 0.09 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.333 0.243 ;

	END

END AOI21x1_ASAP7_75t_L

MACRO AOI21xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI21xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.107 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END AOI21xp33_ASAP7_75t_L

MACRO AOI21xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI21xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.142 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.034 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END AOI21xp5_ASAP7_75t_L

MACRO AOI221x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI221x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.634 0.189 0.738 0.207 ;
			RECT 0.72 0.045 0.738 0.207 ;
			RECT 0.256 0.045 0.738 0.063 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.153 0.217 0.171 ;
			RECT 0.18 0.027 0.198 0.171 ;
			RECT 0.161 0.027 0.198 0.045 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.126 0.149 0.144 ;
			RECT 0.053 0.153 0.09 0.171 ;
			RECT 0.072 0.027 0.09 0.171 ;
			RECT 0.053 0.027 0.09 0.045 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.081 0.325 0.099 ;
			RECT 0.269 0.153 0.306 0.171 ;
			RECT 0.288 0.081 0.306 0.171 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.153 0.487 0.171 ;
			RECT 0.45 0.081 0.468 0.171 ;
			RECT 0.391 0.126 0.468 0.144 ;
			RECT 0.431 0.081 0.468 0.099 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.126 0.636 0.144 ;
			RECT 0.539 0.189 0.576 0.207 ;
			RECT 0.558 0.081 0.576 0.207 ;
			RECT 0.539 0.081 0.576 0.099 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.225 0.716 0.243 ;
			RECT 0.04 0.189 0.5 0.207 ;

	END

END AOI221x1_ASAP7_75t_L

MACRO AOI221xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI221xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.23 0.045 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.201 0.189 0.339 0.207 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AOI221xp5_ASAP7_75t_L

MACRO AOI222xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI222xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.399 0.045 ;
			RECT 0.018 0.189 0.122 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.034 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.342 0.225 0.468 0.243 ;
			RECT 0.342 0.189 0.36 0.243 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI222xp33_ASAP7_75t_L

MACRO AOI22x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI22x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.309 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.038 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.153 0.379 0.171 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.431 0.153 0.468 0.171 ;
			RECT 0.45 0.063 0.468 0.171 ;
			RECT 0.288 0.063 0.468 0.081 ;
			RECT 0.288 0.063 0.306 0.152 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.161 0.189 0.198 0.207 ;
			RECT 0.18 0.099 0.198 0.207 ;
			RECT 0.161 0.099 0.198 0.117 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.252 0.154 ;
			RECT 0.072 0.063 0.252 0.081 ;
			RECT 0.072 0.189 0.109 0.207 ;
			RECT 0.072 0.063 0.09 0.207 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.5 0.243 ;

	END

END AOI22x1_ASAP7_75t_L

MACRO AOI22xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI22xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI22xp33_ASAP7_75t_L

MACRO AOI22xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI22xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.07 0.144 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI22xp5_ASAP7_75t_L

MACRO AOI311xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI311xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.198 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.234 0.243 ;

	END

END AOI311xp33_ASAP7_75t_L

MACRO AOI31xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI31xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.201 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.093 0.225 0.23 0.243 ;

	END

END AOI31xp33_ASAP7_75t_L

MACRO AOI31xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI31xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.585 0.225 0.663 0.243 ;
			RECT 0.585 0.189 0.603 0.243 ;
			RECT 0.202 0.189 0.603 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.202 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.666 0.07 0.684 0.2 ;
			RECT 0.553 0.126 0.684 0.144 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.126 0.419 0.144 ;
			RECT 0.288 0.063 0.325 0.081 ;
			RECT 0.288 0.063 0.306 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.059 0.207 ;
			RECT 0.018 0.027 0.059 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.027 0.663 0.045 ;
			RECT 0.364 0.081 0.608 0.099 ;
			RECT 0.04 0.225 0.554 0.243 ;
			RECT 0.094 0.027 0.447 0.045 ;

	END

END AOI31xp67_ASAP7_75t_L

MACRO AOI321xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI321xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.198 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.225 0.396 0.243 ;
			RECT 0.094 0.189 0.23 0.207 ;

	END

END AOI321xp33_ASAP7_75t_L

MACRO AOI322xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI322xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.189 0.468 0.207 ;
			RECT 0.45 0.027 0.468 0.207 ;
			RECT 0.147 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.165 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.165 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.225 0.45 0.243 ;
			RECT 0.039 0.189 0.284 0.207 ;

	END

END AOI322xp5_ASAP7_75t_L

MACRO AOI32xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI32xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.04 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.058 0.243 ;
			RECT 0.018 0.063 0.058 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.104 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.104 0.063 0.144 0.081 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.222 0.207 ;
			RECT 0.18 0.07 0.198 0.207 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END AOI32xp33_ASAP7_75t_L

MACRO AOI331xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI331xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.417 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.201 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.189 0.393 0.207 ;
			RECT 0.092 0.225 0.339 0.243 ;

	END

END AOI331xp33_ASAP7_75t_L

MACRO AOI332xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI332xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.417 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.201 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.225 0.502 0.243 ;
			RECT 0.092 0.189 0.339 0.207 ;

	END

END AOI332xp33_ASAP7_75t_L

MACRO AOI333xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI333xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.413 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.201 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.225 0.515 0.243 ;
			RECT 0.094 0.189 0.34 0.207 ;

	END

END AOI333xp33_ASAP7_75t_L

MACRO AOI33xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN AOI33xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.201 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.338 0.243 ;

	END

END AOI33xp33_ASAP7_75t_L

MACRO BUFx10_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx10_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.199 0.027 0.738 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.689 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx10_ASAP7_75t_L

MACRO BUFx12_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx12_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.199 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.8 0.144 ;
			RECT 0.094 0.027 0.144 0.045 ;

	END

END BUFx12_ASAP7_75t_L

MACRO BUFx12f_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx12f_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.972 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.31 0.027 0.954 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.074 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.972 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.972 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.243 ;
			RECT 0.261 0.126 0.311 0.144 ;
			RECT 0.094 0.027 0.279 0.045 ;

	END

END BUFx12f_ASAP7_75t_L

MACRO BUFx16f_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx16f_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 1.17 0.243 ;
			RECT 1.152 0.027 1.17 0.243 ;
			RECT 0.31 0.027 1.17 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.06 0.243 ;
			RECT 0.018 0.027 0.06 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.234 0.126 1.124 0.144 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END BUFx16f_ASAP7_75t_L

MACRO BUFx24_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx24_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.62 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 1.602 0.243 ;
			RECT 1.584 0.027 1.602 0.243 ;
			RECT 0.31 0.027 1.602 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.62 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.62 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.234 0.126 1.553 0.144 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END BUFx24_ASAP7_75t_L

MACRO BUFx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.145 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.203 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx2_ASAP7_75t_L

MACRO BUFx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.145 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.26 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx3_ASAP7_75t_L

MACRO BUFx4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.357 0.243 ;
			RECT 0.339 0.027 0.357 0.243 ;
			RECT 0.145 0.027 0.357 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.314 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx4_ASAP7_75t_L

MACRO BUFx4f_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx4f_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.199 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.098 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.367 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx4f_ASAP7_75t_L

MACRO BUFx5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.145 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.368 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx5_ASAP7_75t_L

MACRO BUFx6f_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx6f_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.202 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.473 0.144 ;
			RECT 0.094 0.027 0.144 0.045 ;

	END

END BUFx6f_ASAP7_75t_L

MACRO BUFx8_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN BUFx8_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.202 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.098 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.581 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx8_ASAP7_75t_L

MACRO CKINVDCx10_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx10_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.296 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.224 0.243 ;
			RECT 1.206 0.063 1.224 0.243 ;
			RECT 1.174 0.063 1.224 0.081 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.17 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.296 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.296 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx10_ASAP7_75t_L

MACRO CKINVDCx11_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx11_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.31 0.243 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.354 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx11_ASAP7_75t_L

MACRO CKINVDCx12_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx12_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.31 0.243 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.354 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx12_ASAP7_75t_L

MACRO CKINVDCx14_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx14_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.512 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.44 0.243 ;
			RECT 1.422 0.063 1.44 0.243 ;
			RECT 1.39 0.063 1.44 0.081 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.397 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.512 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.512 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx14_ASAP7_75t_L

MACRO CKINVDCx16_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx16_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.62 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 1.548 0.243 ;
			RECT 1.53 0.063 1.548 0.243 ;
			RECT 1.498 0.063 1.548 0.081 ;
			RECT 1.368 0.063 1.418 0.081 ;
			RECT 1.368 0.063 1.386 0.243 ;
			RECT 1.098 0.063 1.116 0.243 ;
			RECT 1.066 0.063 1.116 0.081 ;
			RECT 0.936 0.063 0.986 0.081 ;
			RECT 0.936 0.063 0.954 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.634 0.063 0.684 0.081 ;
			RECT 0.504 0.063 0.554 0.081 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.202 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.122 0.081 ;
			RECT 0.072 0.063 0.09 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.412 0.126 1.505 0.144 ;
			RECT 1.444 0.027 1.462 0.144 ;
			RECT 0.158 0.027 1.462 0.045 ;
			RECT 0.98 0.126 1.072 0.144 ;
			RECT 1.017 0.027 1.035 0.144 ;
			RECT 0.547 0.126 0.639 0.144 ;
			RECT 0.584 0.027 0.602 0.144 ;
			RECT 0.126 0.126 0.208 0.144 ;
			RECT 0.158 0.027 0.176 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.62 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.62 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.26 0.126 1.316 0.144 ;
			RECT 1.26 0.09 1.278 0.144 ;
			RECT 1.174 0.09 1.326 0.108 ;
			RECT 1.155 0.162 1.31 0.18 ;
			RECT 1.206 0.126 1.224 0.18 ;
			RECT 1.166 0.126 1.224 0.144 ;
			RECT 0.742 0.162 0.897 0.18 ;
			RECT 0.828 0.126 0.846 0.18 ;
			RECT 0.828 0.126 0.886 0.144 ;
			RECT 0.736 0.126 0.792 0.144 ;
			RECT 0.774 0.09 0.792 0.144 ;
			RECT 0.726 0.09 0.878 0.108 ;
			RECT 0.31 0.162 0.465 0.18 ;
			RECT 0.396 0.126 0.414 0.18 ;
			RECT 0.396 0.126 0.454 0.144 ;
			RECT 0.304 0.126 0.36 0.144 ;
			RECT 0.342 0.09 0.36 0.144 ;
			RECT 0.294 0.09 0.446 0.108 ;

	END

END CKINVDCx16_ASAP7_75t_L

MACRO CKINVDCx20_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx20_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.052 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 1.98 0.243 ;
			RECT 1.962 0.063 1.98 0.243 ;
			RECT 1.93 0.063 1.98 0.081 ;
			RECT 1.8 0.063 1.85 0.081 ;
			RECT 1.8 0.063 1.818 0.243 ;
			RECT 1.53 0.063 1.548 0.243 ;
			RECT 1.498 0.063 1.548 0.081 ;
			RECT 1.368 0.063 1.418 0.081 ;
			RECT 1.368 0.063 1.386 0.243 ;
			RECT 1.098 0.063 1.116 0.243 ;
			RECT 1.066 0.063 1.116 0.081 ;
			RECT 0.936 0.063 0.986 0.081 ;
			RECT 0.936 0.063 0.954 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.634 0.063 0.684 0.081 ;
			RECT 0.504 0.063 0.554 0.081 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.202 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.122 0.081 ;
			RECT 0.072 0.063 0.09 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.844 0.126 1.937 0.144 ;
			RECT 1.876 0.027 1.894 0.144 ;
			RECT 0.158 0.027 1.894 0.045 ;
			RECT 1.412 0.126 1.505 0.144 ;
			RECT 1.444 0.027 1.462 0.144 ;
			RECT 0.98 0.126 1.072 0.144 ;
			RECT 1.017 0.027 1.035 0.144 ;
			RECT 0.547 0.126 0.639 0.144 ;
			RECT 0.584 0.027 0.602 0.144 ;
			RECT 0.126 0.126 0.208 0.144 ;
			RECT 0.158 0.027 0.176 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.052 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.052 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.692 0.126 1.748 0.144 ;
			RECT 1.692 0.09 1.71 0.144 ;
			RECT 1.606 0.09 1.758 0.108 ;
			RECT 1.587 0.162 1.742 0.18 ;
			RECT 1.638 0.126 1.656 0.18 ;
			RECT 1.598 0.126 1.656 0.144 ;
			RECT 1.26 0.126 1.316 0.144 ;
			RECT 1.26 0.09 1.278 0.144 ;
			RECT 1.174 0.09 1.326 0.108 ;
			RECT 1.155 0.162 1.31 0.18 ;
			RECT 1.206 0.126 1.224 0.18 ;
			RECT 1.166 0.126 1.224 0.144 ;
			RECT 0.742 0.162 0.897 0.18 ;
			RECT 0.828 0.126 0.846 0.18 ;
			RECT 0.828 0.126 0.886 0.144 ;
			RECT 0.736 0.126 0.792 0.144 ;
			RECT 0.774 0.09 0.792 0.144 ;
			RECT 0.726 0.09 0.878 0.108 ;
			RECT 0.31 0.162 0.465 0.18 ;
			RECT 0.396 0.126 0.414 0.18 ;
			RECT 0.396 0.126 0.454 0.144 ;
			RECT 0.304 0.126 0.36 0.144 ;
			RECT 0.342 0.09 0.36 0.144 ;
			RECT 0.294 0.09 0.446 0.108 ;

	END

END CKINVDCx20_ASAP7_75t_L

MACRO CKINVDCx5p33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx5p33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.094 0.243 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.138 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx5p33_ASAP7_75t_L

MACRO CKINVDCx6p67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx6p67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.296 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.224 0.243 ;
			RECT 1.206 0.063 1.224 0.243 ;
			RECT 1.174 0.063 1.224 0.081 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.17 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.296 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.296 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx6p67_ASAP7_75t_L

MACRO CKINVDCx8_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx8_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.094 0.243 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.138 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx8_ASAP7_75t_L

MACRO CKINVDCx9p33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN CKINVDCx9p33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.512 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.44 0.243 ;
			RECT 1.422 0.063 1.44 0.243 ;
			RECT 1.39 0.063 1.44 0.081 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.397 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.512 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.512 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx9p33_ASAP7_75t_L

MACRO DECAPx10_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN DECAPx10_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.558 0.045 0.576 0.15 ;
			RECT 0.558 0.045 1.148 0.063 ;
			RECT 0.04 0.207 0.63 0.225 ;
			RECT 0.612 0.121 0.63 0.225 ;

	END

END DECAPx10_ASAP7_75t_L

MACRO DECAPx1_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN DECAPx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.207 0.144 0.225 ;
			RECT 0.126 0.121 0.144 0.225 ;
			RECT 0.072 0.045 0.09 0.15 ;
			RECT 0.072 0.045 0.122 0.063 ;

	END

END DECAPx1_ASAP7_75t_L

MACRO DECAPx2_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN DECAPx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.045 0.144 0.15 ;
			RECT 0.126 0.045 0.284 0.063 ;
			RECT 0.04 0.207 0.198 0.225 ;
			RECT 0.18 0.121 0.198 0.225 ;

	END

END DECAPx2_ASAP7_75t_L

MACRO DECAPx2b_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN DECAPx2b_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.162 0.249 0.18 ;
			RECT 0.18 0.126 0.198 0.18 ;
			RECT 0.18 0.126 0.238 0.144 ;
			RECT 0.088 0.126 0.144 0.144 ;
			RECT 0.126 0.09 0.144 0.144 ;
			RECT 0.078 0.09 0.23 0.108 ;

	END

END DECAPx2b_ASAP7_75t_L

MACRO DECAPx4_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN DECAPx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.234 0.045 0.252 0.15 ;
			RECT 0.234 0.045 0.5 0.063 ;
			RECT 0.04 0.207 0.306 0.225 ;
			RECT 0.288 0.121 0.306 0.225 ;

	END

END DECAPx4_ASAP7_75t_L

MACRO DECAPx6_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN DECAPx6_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.342 0.045 0.36 0.15 ;
			RECT 0.342 0.045 0.716 0.063 ;
			RECT 0.04 0.207 0.414 0.225 ;
			RECT 0.396 0.121 0.414 0.225 ;

	END

END DECAPx6_ASAP7_75t_L

MACRO DFFASRHQNx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFASRHQNx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.336 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.336 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.182 0.117 0.236 ;
			RECT 0.072 0.182 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN RESETN
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.632 0.144 1.067 0.162 ;
			LAYER M1 ;
			RECT 1.044 0.102 1.062 0.167 ;
			RECT 0.612 0.072 0.668 0.09 ;
			RECT 0.612 0.144 0.662 0.162 ;
			RECT 0.612 0.072 0.63 0.162 ;
			LAYER V1 ;
			RECT 0.637 0.144 0.655 0.162 ;
			RECT 1.044 0.144 1.062 0.162 ;

		END 

	END RESETN
	PIN SETN
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.783 0.18 1.067 0.198 ;
			LAYER M1 ;
			RECT 0.774 0.18 0.811 0.198 ;
			RECT 0.774 0.097 0.792 0.198 ;
			LAYER V1 ;
			RECT 0.788 0.18 0.806 0.198 ;

		END 

	END SETN
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.963 0.036 0.981 0.234 ;
			RECT 0.963 0.036 1.008 0.054 ;
			RECT 0.855 0.222 0.936 0.24 ;
			RECT 0.918 0.053 0.936 0.24 ;
			RECT 0.693 0.036 0.711 0.212 ;
			RECT 0.558 0.036 0.576 0.106 ;
			RECT 0.558 0.036 0.77 0.054 ;
			RECT 0.486 0.18 0.547 0.198 ;
			RECT 0.486 0.027 0.504 0.198 ;
			RECT 0.418 0.027 0.504 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.142 0.027 0.198 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.018 0.108 0.047 0.126 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 1.314 0.103 1.332 0.18 ;
			RECT 1.17 0.216 1.202 0.234 ;
			RECT 1.098 0.102 1.116 0.167 ;
			RECT 0.882 0.067 0.9 0.173 ;
			RECT 0.829 0.103 0.847 0.171 ;
			RECT 0.778 0.216 0.819 0.234 ;
			RECT 0.729 0.137 0.747 0.203 ;
			RECT 0.415 0.225 0.608 0.243 ;
			RECT 0.45 0.103 0.468 0.151 ;
			RECT 0.396 0.067 0.414 0.15 ;
			RECT 0.369 0.169 0.387 0.216 ;
			RECT 0.342 0.103 0.36 0.15 ;
			RECT 0.142 0.07 0.16 0.164 ;
			LAYER M2 ;
			RECT 0.913 0.108 1.337 0.126 ;
			RECT 0.783 0.216 1.198 0.234 ;
			RECT 0.741 0.036 1.008 0.054 ;
			RECT 0.018 0.072 0.926 0.09 ;
			RECT 0.175 0.108 0.852 0.126 ;
			RECT 0.364 0.18 0.752 0.198 ;
			LAYER V1 ;
			RECT 1.314 0.108 1.332 0.126 ;
			RECT 1.175 0.216 1.193 0.234 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 0.985 0.036 1.003 0.054 ;
			RECT 0.918 0.108 0.936 0.126 ;
			RECT 0.882 0.072 0.9 0.09 ;
			RECT 0.829 0.108 0.847 0.126 ;
			RECT 0.788 0.216 0.806 0.234 ;
			RECT 0.746 0.036 0.764 0.054 ;
			RECT 0.729 0.18 0.747 0.198 ;
			RECT 0.512 0.18 0.53 0.198 ;
			RECT 0.45 0.108 0.468 0.126 ;
			RECT 0.396 0.072 0.414 0.09 ;
			RECT 0.369 0.18 0.387 0.198 ;
			RECT 0.342 0.108 0.36 0.126 ;
			RECT 0.18 0.108 0.198 0.126 ;
			RECT 0.142 0.072 0.16 0.09 ;
			RECT 0.018 0.072 0.036 0.09 ;

	END

END DFFASRHQNx1_ASAP7_75t_L

MACRO DFFHQNx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFHQNx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 1.012 0.027 1.062 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx1_ASAP7_75t_L

MACRO DFFHQNx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFHQNx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.216 1.117 0.234 ;
			RECT 1.099 0.036 1.117 0.234 ;
			RECT 1.012 0.036 1.117 0.054 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx2_ASAP7_75t_L

MACRO DFFHQNx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFHQNx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.171 0.243 ;
			RECT 1.153 0.027 1.171 0.243 ;
			RECT 1.012 0.027 1.171 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx3_ASAP7_75t_L

MACRO DFFHQx4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFHQx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.125 0.225 1.333 0.243 ;
			RECT 1.313 0.027 1.333 0.243 ;
			RECT 1.125 0.027 1.333 0.045 ;
			RECT 1.125 0.201 1.143 0.243 ;
			RECT 1.125 0.027 1.143 0.069 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.012 0.225 1.098 0.243 ;
			RECT 1.08 0.027 1.098 0.243 ;
			RECT 1.08 0.127 1.175 0.145 ;
			RECT 1.012 0.027 1.098 0.045 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQx4_ASAP7_75t_L

MACRO DFFLQNx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFLQNx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 1.012 0.027 1.062 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx1_ASAP7_75t_L

MACRO DFFLQNx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFLQNx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.115 0.243 ;
			RECT 1.097 0.027 1.115 0.243 ;
			RECT 1.012 0.027 1.115 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx2_ASAP7_75t_L

MACRO DFFLQNx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFLQNx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.171 0.243 ;
			RECT 1.153 0.027 1.171 0.243 ;
			RECT 1.011 0.027 1.171 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx3_ASAP7_75t_L

MACRO DFFLQx4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DFFLQx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.125 0.225 1.333 0.243 ;
			RECT 1.313 0.027 1.333 0.243 ;
			RECT 1.125 0.027 1.333 0.045 ;
			RECT 1.125 0.201 1.143 0.243 ;
			RECT 1.125 0.027 1.143 0.069 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.012 0.225 1.098 0.243 ;
			RECT 1.08 0.027 1.098 0.243 ;
			RECT 1.08 0.127 1.175 0.145 ;
			RECT 1.012 0.027 1.098 0.045 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQx4_ASAP7_75t_L

MACRO DHLx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DHLx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.742 0.027 0.792 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.72 0.122 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.743 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx1_ASAP7_75t_L

MACRO DHLx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DHLx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.741 0.216 0.85 0.234 ;
			RECT 0.832 0.036 0.85 0.234 ;
			RECT 0.742 0.036 0.85 0.054 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.72 0.09 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.797 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx2_ASAP7_75t_L

MACRO DHLx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DHLx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.918 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.688 0.225 0.9 0.243 ;
			RECT 0.882 0.027 0.9 0.243 ;
			RECT 0.688 0.027 0.9 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.918 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.918 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.828 0.09 0.846 0.167 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.72 0.09 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.851 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx3_ASAP7_75t_L

MACRO DLLx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DLLx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.735 0.027 0.792 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.72 0.106 0.738 0.2 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.743 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx1_ASAP7_75t_L

MACRO DLLx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DLLx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.688 0.225 0.847 0.243 ;
			RECT 0.829 0.027 0.847 0.243 ;
			RECT 0.688 0.027 0.847 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.8 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx2_ASAP7_75t_L

MACRO DLLx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN DLLx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.918 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.216 0.901 0.234 ;
			RECT 0.882 0.036 0.901 0.234 ;
			RECT 0.742 0.036 0.901 0.054 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.918 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.918 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.8 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx3_ASAP7_75t_L

MACRO FAx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN FAx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN CON
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.128 0.072 0.543 0.09 ;
			LAYER M1 ;
			RECT 0.515 0.072 0.543 0.09 ;
			RECT 0.504 0.09 0.533 0.108 ;
			RECT 0.504 0.09 0.522 0.149 ;
			RECT 0.124 0.072 0.282 0.09 ;
			RECT 0.124 0.189 0.23 0.207 ;
			RECT 0.124 0.072 0.142 0.207 ;
			LAYER V1 ;
			RECT 0.133 0.072 0.151 0.09 ;
			RECT 0.52 0.072 0.538 0.09 ;

		END 

	END CON
	PIN SN
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.324 0.225 0.495 0.243 ;
			RECT 0.477 0.184 0.495 0.243 ;
			RECT 0.477 0.027 0.495 0.068 ;
			RECT 0.324 0.027 0.495 0.045 ;
			RECT 0.324 0.027 0.342 0.243 ;

		END 

	END SN
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.059 0.18 0.627 0.198 ;
			LAYER M1 ;
			RECT 0.599 0.18 0.63 0.198 ;
			RECT 0.612 0.121 0.63 0.198 ;
			RECT 0.383 0.18 0.414 0.198 ;
			RECT 0.396 0.121 0.414 0.198 ;
			RECT 0.059 0.18 0.09 0.198 ;
			RECT 0.072 0.121 0.09 0.198 ;
			LAYER V1 ;
			RECT 0.064 0.18 0.082 0.198 ;
			RECT 0.388 0.18 0.406 0.198 ;
			RECT 0.604 0.18 0.622 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.167 0.144 0.689 0.162 ;
			LAYER M1 ;
			RECT 0.666 0.121 0.684 0.167 ;
			RECT 0.288 0.121 0.306 0.167 ;
			RECT 0.167 0.144 0.198 0.162 ;
			RECT 0.18 0.121 0.198 0.162 ;
			LAYER V1 ;
			RECT 0.172 0.144 0.19 0.162 ;
			RECT 0.288 0.144 0.306 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;

		END 

	END B
	PIN CI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.108 0.587 0.126 ;
			LAYER M1 ;
			RECT 0.558 0.108 0.587 0.126 ;
			RECT 0.558 0.108 0.576 0.149 ;
			RECT 0.45 0.103 0.468 0.149 ;
			RECT 0.226 0.108 0.263 0.126 ;
			RECT 0.234 0.108 0.252 0.149 ;
			LAYER V1 ;
			RECT 0.234 0.108 0.252 0.126 ;
			RECT 0.45 0.108 0.468 0.126 ;
			RECT 0.564 0.108 0.582 0.126 ;

		END 

	END CI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.027 0.662 0.045 ;
			RECT 0.526 0.225 0.662 0.243 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END FAx1_ASAP7_75t_L

MACRO FILLER_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN FILLER_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.108 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.108 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.108 0.279 ;

		END 

	END VDD

END FILLER_ASAP7_75t_L

MACRO FILLERxp5_ASAP7_75t_L
	CLASS CORE SPACER ;
	FOREIGN FILLERxp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.054 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.054 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.054 0.279 ;

		END 

	END VDD

END FILLERxp5_ASAP7_75t_L

MACRO HAxp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN HAxp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN CON
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.162 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.075 0.18 0.243 ;

		END 

	END CON
	PIN SN
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.423 0.027 0.468 0.045 ;

		END 

	END SN
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.15 ;
			RECT 0.207 0.063 0.36 0.081 ;
			RECT 0.207 0.027 0.225 0.081 ;
			RECT 0.018 0.027 0.225 0.045 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.027 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.106 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.387 0.045 ;

	END

END HAxp5_ASAP7_75t_L

MACRO HB1xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN HB1xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.117 0.243 ;
			RECT 0.099 0.153 0.117 0.243 ;
			RECT 0.099 0.153 0.144 0.171 ;
			RECT 0.126 0.099 0.144 0.171 ;
			RECT 0.099 0.099 0.144 0.117 ;
			RECT 0.099 0.027 0.117 0.117 ;
			RECT 0.04 0.027 0.117 0.045 ;

	END

END HB1xp67_ASAP7_75t_L

MACRO HB2xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN HB2xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.202 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.04 0.027 0.144 0.045 ;

	END

END HB2xp67_ASAP7_75t_L

MACRO HB3xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN HB3xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.256 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.18 0.126 0.257 0.144 ;
			RECT 0.04 0.027 0.198 0.045 ;

	END

END HB3xp67_ASAP7_75t_L

MACRO HB4xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN HB4xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.081 0.055 0.099 ;
			RECT 0.018 0.081 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.18 0.126 0.311 0.144 ;
			RECT 0.04 0.027 0.198 0.045 ;

	END

END HB4xp67_ASAP7_75t_L

MACRO ICGx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.972 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.879 0.027 0.954 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.972 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.972 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx1_ASAP7_75t_L

MACRO ICGx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.026 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 1.008 0.243 ;
			RECT 0.99 0.027 1.008 0.243 ;
			RECT 0.879 0.027 1.008 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.026 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.026 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx2_ASAP7_75t_L

MACRO ICGx2p67DC_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx2p67DC_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx2p67DC_ASAP7_75t_L

MACRO ICGx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.879 0.027 1.062 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx3_ASAP7_75t_L

MACRO ICGx4DC_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx4DC_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx4DC_ASAP7_75t_L

MACRO ICGx4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.89 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.889 0.027 1.062 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx4_ASAP7_75t_L

MACRO ICGx5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.89 0.225 1.17 0.243 ;
			RECT 1.152 0.027 1.17 0.243 ;
			RECT 0.889 0.027 1.17 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx5_ASAP7_75t_L

MACRO ICGx5p33DC_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx5p33DC_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx5p33DC_ASAP7_75t_L

MACRO ICGx6p67DC_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx6p67DC_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx6p67DC_ASAP7_75t_L

MACRO ICGx8DC_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN ICGx8DC_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx8DC_ASAP7_75t_L

MACRO INVx11_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx11_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.094 0.027 0.684 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD

END INVx11_ASAP7_75t_L

MACRO INVx13_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx13_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.094 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD

END INVx13_ASAP7_75t_L

MACRO INVx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVx1_ASAP7_75t_L

MACRO INVx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END INVx2_ASAP7_75t_L

MACRO INVx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.094 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END INVx3_ASAP7_75t_L

MACRO INVx4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END INVx4_ASAP7_75t_L

MACRO INVx5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.094 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END INVx5_ASAP7_75t_L

MACRO INVx6_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx6_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.094 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD

END INVx6_ASAP7_75t_L

MACRO INVx8_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVx8_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.094 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD

END INVx8_ASAP7_75t_L

MACRO INVxp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVxp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVxp33_ASAP7_75t_L

MACRO INVxp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN INVxp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVxp67_ASAP7_75t_L

MACRO MAJIxp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN MAJIxp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.255 0.189 0.361 0.207 ;
			RECT 0.343 0.063 0.361 0.207 ;
			RECT 0.255 0.063 0.361 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.126 0.257 0.144 ;
			RECT 0.018 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.027 0.338 0.045 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END MAJIxp5_ASAP7_75t_L

MACRO MAJx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN MAJx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.364 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.333 0.207 ;
			RECT 0.315 0.106 0.333 0.207 ;
			RECT 0.283 0.126 0.333 0.144 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.121 0.126 0.198 0.144 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.063 0.036 0.207 ;
			RECT 0.368 0.063 0.386 0.149 ;
			RECT 0.018 0.063 0.386 0.081 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END MAJx2_ASAP7_75t_L

MACRO MAJx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN MAJx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.504 0.243 ;
			RECT 0.364 0.027 0.504 0.045 ;
			RECT 0.45 0.027 0.468 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.333 0.207 ;
			RECT 0.315 0.106 0.333 0.207 ;
			RECT 0.283 0.126 0.333 0.144 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.121 0.126 0.198 0.144 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.063 0.036 0.207 ;
			RECT 0.368 0.063 0.386 0.149 ;
			RECT 0.018 0.063 0.386 0.081 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END MAJx3_ASAP7_75t_L

MACRO NAND2x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND2x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.202 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.065 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END NAND2x1_ASAP7_75t_L

MACRO NAND2x1p5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND2x1p5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.261 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.063 0.338 0.081 ;
			RECT 0.094 0.027 0.225 0.045 ;

	END

END NAND2x1p5_ASAP7_75t_L

MACRO NAND2x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND2x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.418 0.063 0.522 0.081 ;
			RECT 0.018 0.063 0.122 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.242 0.189 0.279 0.207 ;
			RECT 0.261 0.106 0.279 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.177 ;
			RECT 0.322 0.099 0.468 0.117 ;
			RECT 0.322 0.063 0.34 0.117 ;
			RECT 0.2 0.063 0.34 0.081 ;
			RECT 0.072 0.099 0.218 0.117 ;
			RECT 0.2 0.063 0.218 0.117 ;
			RECT 0.072 0.189 0.109 0.207 ;
			RECT 0.072 0.099 0.09 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.5 0.045 ;

	END

END NAND2x2_ASAP7_75t_L

MACRO NAND2xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND2xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.143 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NAND2xp33_ASAP7_75t_L

MACRO NAND2xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND2xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.143 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.106 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NAND2xp5_ASAP7_75t_L

MACRO NAND2xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND2xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.202 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.106 0.252 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END NAND2xp67_ASAP7_75t_L

MACRO NAND3x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND3x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.418 0.063 0.576 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.402 0.18 0.468 0.198 ;
			RECT 0.45 0.108 0.468 0.198 ;
			RECT 0.4 0.108 0.468 0.126 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.243 0.18 0.306 0.198 ;
			RECT 0.288 0.108 0.306 0.198 ;
			RECT 0.246 0.108 0.306 0.126 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.061 0.103 0.079 0.203 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.5 0.045 ;
			RECT 0.094 0.063 0.338 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END NAND3x1_ASAP7_75t_L

MACRO NAND3x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND3x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 1.062 0.243 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.904 0.063 1.062 0.081 ;
			RECT 0.018 0.063 0.176 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.169 0.18 0.908 0.198 ;
			LAYER M1 ;
			RECT 0.866 0.189 0.903 0.207 ;
			RECT 0.885 0.108 0.903 0.207 ;
			RECT 0.174 0.189 0.211 0.207 ;
			RECT 0.174 0.106 0.192 0.207 ;
			LAYER V1 ;
			RECT 0.174 0.18 0.192 0.198 ;
			RECT 0.885 0.18 0.903 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.338 0.189 0.743 0.207 ;
			RECT 0.725 0.106 0.743 0.207 ;
			RECT 0.338 0.106 0.356 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.547 0.106 0.565 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.742 0.027 0.986 0.045 ;
			RECT 0.256 0.063 0.824 0.081 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.094 0.027 0.338 0.045 ;

	END

END NAND3x2_ASAP7_75t_L

MACRO NAND3xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND3xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END NAND3xp33_ASAP7_75t_L

MACRO NAND4xp25_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND4xp25_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.256 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END NAND4xp25_ASAP7_75t_L

MACRO NAND4xp75_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND4xp75_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.738 0.243 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.58 0.063 0.738 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.106 0.63 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.101 0.549 0.119 ;
			RECT 0.531 0.07 0.549 0.119 ;
			RECT 0.504 0.101 0.522 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.101 0.306 0.2 ;
			RECT 0.207 0.101 0.306 0.119 ;
			RECT 0.207 0.07 0.225 0.119 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.057 0.243 ;
			RECT 0.018 0.027 0.057 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.412 0.027 0.666 0.045 ;
			RECT 0.256 0.063 0.499 0.081 ;
			RECT 0.092 0.027 0.34 0.045 ;

	END

END NAND4xp75_ASAP7_75t_L

MACRO NAND5xp2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NAND5xp2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.009 0.225 0.317 0.243 ;
			RECT 0.009 0.027 0.07 0.045 ;
			RECT 0.009 0.027 0.027 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.2 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END NAND5xp2_ASAP7_75t_L

MACRO NOR2x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR2x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.23 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END NOR2x1_ASAP7_75t_L

MACRO NOR2x1p5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR2x1p5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.094 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.063 0.163 0.081 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.338 0.207 ;
			RECT 0.094 0.225 0.225 0.243 ;

	END

END NOR2x1p5_ASAP7_75t_L

MACRO NOR2x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR2x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.018 0.027 0.522 0.045 ;
			RECT 0.018 0.189 0.122 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.063 0.279 0.164 ;
			RECT 0.242 0.063 0.279 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.322 0.153 0.468 0.171 ;
			RECT 0.45 0.093 0.468 0.171 ;
			RECT 0.2 0.189 0.34 0.207 ;
			RECT 0.322 0.153 0.34 0.207 ;
			RECT 0.2 0.153 0.218 0.207 ;
			RECT 0.072 0.153 0.218 0.171 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.5 0.243 ;

	END

END NOR2x2_ASAP7_75t_L

MACRO NOR2xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR2xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.143 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.094 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NOR2xp33_ASAP7_75t_L

MACRO NOR2xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR2xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.127 0.095 0.145 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.063 0.163 0.081 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END NOR2xp67_ASAP7_75t_L

MACRO NOR3x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR3x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.202 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.153 0.468 0.171 ;
			RECT 0.45 0.063 0.468 0.171 ;
			RECT 0.396 0.063 0.468 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.153 0.306 0.171 ;
			RECT 0.288 0.063 0.306 0.171 ;
			RECT 0.234 0.063 0.306 0.081 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.225 0.5 0.243 ;
			RECT 0.094 0.189 0.338 0.207 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END NOR3x1_ASAP7_75t_L

MACRO NOR3x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR3x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.904 0.189 1.062 0.207 ;
			RECT 1.044 0.027 1.062 0.207 ;
			RECT 0.018 0.027 1.062 0.045 ;
			RECT 0.018 0.189 0.176 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.169 0.072 0.908 0.09 ;
			LAYER M1 ;
			RECT 0.885 0.063 0.903 0.162 ;
			RECT 0.866 0.063 0.903 0.081 ;
			RECT 0.174 0.063 0.211 0.081 ;
			RECT 0.174 0.063 0.192 0.164 ;
			LAYER V1 ;
			RECT 0.174 0.072 0.192 0.09 ;
			RECT 0.885 0.072 0.903 0.09 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.725 0.063 0.743 0.164 ;
			RECT 0.338 0.063 0.743 0.081 ;
			RECT 0.338 0.063 0.356 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.547 0.106 0.565 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.742 0.225 0.986 0.243 ;
			RECT 0.256 0.189 0.824 0.207 ;
			RECT 0.418 0.225 0.662 0.243 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END NOR3x2_ASAP7_75t_L

MACRO NOR3xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR3xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.176 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END NOR3xp33_ASAP7_75t_L

MACRO NOR4xp25_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR4xp25_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.04 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END NOR4xp25_ASAP7_75t_L

MACRO NOR4xp75_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR4xp75_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.58 0.189 0.738 0.207 ;
			RECT 0.72 0.027 0.738 0.207 ;
			RECT 0.094 0.027 0.738 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.07 0.63 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.531 0.151 0.549 0.2 ;
			RECT 0.504 0.151 0.549 0.169 ;
			RECT 0.504 0.07 0.522 0.169 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.151 0.306 0.169 ;
			RECT 0.288 0.07 0.306 0.169 ;
			RECT 0.207 0.151 0.225 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.057 0.243 ;
			RECT 0.018 0.027 0.057 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.412 0.225 0.666 0.243 ;
			RECT 0.256 0.189 0.499 0.207 ;
			RECT 0.092 0.225 0.34 0.243 ;

	END

END NOR4xp75_ASAP7_75t_L

MACRO NOR5xp2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN NOR5xp2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.017 0.027 0.338 0.045 ;
			RECT 0.017 0.225 0.07 0.243 ;
			RECT 0.017 0.027 0.037 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END NOR5xp2_ASAP7_75t_L

MACRO O2A1O1Ixp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN O2A1O1Ixp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.206 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.225 0.243 ;
			RECT 0.04 0.063 0.176 0.081 ;

	END

END O2A1O1Ixp33_ASAP7_75t_L

MACRO O2A1O1Ixp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN O2A1O1Ixp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.315 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.252 0.164 ;
			RECT 0.072 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.189 0.338 0.207 ;
			RECT 0.148 0.027 0.279 0.045 ;
			RECT 0.094 0.225 0.23 0.243 ;

	END

END O2A1O1Ixp5_ASAP7_75t_L

MACRO OA211x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA211x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.296 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.286 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.234 0.189 0.306 0.207 ;
			RECT 0.288 0.063 0.306 0.207 ;
			RECT 0.099 0.063 0.306 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OA211x2_ASAP7_75t_L

MACRO OA21x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA21x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.256 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.153 0.239 0.171 ;
			RECT 0.18 0.106 0.198 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.225 0.224 0.243 ;
			RECT 0.206 0.189 0.224 0.243 ;
			RECT 0.206 0.189 0.306 0.207 ;
			RECT 0.288 0.063 0.306 0.207 ;
			RECT 0.099 0.063 0.306 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OA21x2_ASAP7_75t_L

MACRO OA221x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA221x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.225 0.117 0.243 ;
			RECT 0.099 0.189 0.117 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.099 0.252 0.207 ;
			RECT 0.215 0.099 0.252 0.117 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.593 0.189 0.63 0.207 ;
			RECT 0.612 0.099 0.63 0.207 ;
			RECT 0.593 0.099 0.63 0.117 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.099 0.522 0.207 ;
			RECT 0.485 0.099 0.522 0.117 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.72 0.189 0.757 0.207 ;
			RECT 0.72 0.099 0.757 0.117 ;
			RECT 0.72 0.099 0.738 0.207 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.144 0.225 0.846 0.243 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.144 0.126 0.162 0.243 ;
			RECT 0.121 0.126 0.162 0.144 ;
			RECT 0.741 0.063 0.846 0.081 ;
			RECT 0.472 0.027 0.824 0.045 ;
			RECT 0.202 0.063 0.668 0.081 ;

	END

END OA221x2_ASAP7_75t_L

MACRO OA222x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA222x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.531 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.526 0.027 0.63 0.045 ;
			RECT 0.531 0.189 0.549 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.009 0.225 0.504 0.243 ;
			RECT 0.486 0.126 0.504 0.243 ;
			RECT 0.009 0.063 0.027 0.243 ;
			RECT 0.486 0.126 0.554 0.144 ;
			RECT 0.009 0.063 0.122 0.081 ;
			RECT 0.202 0.063 0.36 0.081 ;
			RECT 0.342 0.027 0.36 0.081 ;
			RECT 0.342 0.027 0.468 0.045 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OA222x2_ASAP7_75t_L

MACRO OA22x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA22x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.071 0.225 0.122 0.243 ;
			RECT 0.071 0.027 0.122 0.045 ;
			RECT 0.071 0.027 0.091 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.236 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.063 0.414 0.2 ;
			RECT 0.367 0.063 0.414 0.081 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.18 0.225 0.392 0.243 ;
			RECT 0.18 0.063 0.198 0.243 ;
			RECT 0.137 0.126 0.198 0.144 ;
			RECT 0.18 0.063 0.333 0.081 ;
			RECT 0.256 0.027 0.5 0.045 ;

	END

END OA22x2_ASAP7_75t_L

MACRO OA31x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA31x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.693 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.053 0.189 0.09 0.207 ;
			RECT 0.072 0.099 0.09 0.207 ;
			RECT 0.053 0.099 0.09 0.117 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.126 0.189 0.163 0.207 ;
			RECT 0.126 0.106 0.144 0.207 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.126 0.414 0.144 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.323 0.063 0.36 0.081 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.153 0.522 0.171 ;
			RECT 0.504 0.106 0.522 0.171 ;

		END 

	END B1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.369 0.189 0.576 0.207 ;
			RECT 0.558 0.063 0.576 0.207 ;
			RECT 0.558 0.126 0.667 0.144 ;
			RECT 0.418 0.063 0.576 0.081 ;
			RECT 0.317 0.225 0.446 0.243 ;
			RECT 0.317 0.189 0.335 0.243 ;
			RECT 0.202 0.189 0.335 0.207 ;
			RECT 0.094 0.027 0.5 0.045 ;
			RECT 0.04 0.063 0.284 0.081 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END OA31x2_ASAP7_75t_L

MACRO OA331x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA331x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.166 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.099 0.186 0.117 0.243 ;
			RECT 0.072 0.186 0.117 0.204 ;
			RECT 0.072 0.115 0.09 0.204 ;
			RECT 0.471 0.063 0.522 0.081 ;
			RECT 0.234 0.063 0.393 0.081 ;
			RECT 0.234 0.027 0.252 0.081 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.308 0.027 0.447 0.045 ;

	END

END OA331x1_ASAP7_75t_L

MACRO OA331x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA331x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.045 0.225 0.122 0.243 ;
			RECT 0.045 0.027 0.122 0.045 ;
			RECT 0.045 0.027 0.063 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.166 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.153 0.186 0.171 0.243 ;
			RECT 0.126 0.186 0.171 0.204 ;
			RECT 0.126 0.115 0.144 0.204 ;
			RECT 0.525 0.063 0.576 0.081 ;
			RECT 0.288 0.063 0.447 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.202 0.027 0.306 0.045 ;
			RECT 0.362 0.027 0.501 0.045 ;

	END

END OA331x2_ASAP7_75t_L

MACRO OA332x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA332x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.094 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.126 0.189 0.144 0.243 ;
			RECT 0.072 0.189 0.144 0.207 ;
			RECT 0.072 0.119 0.09 0.207 ;
			RECT 0.471 0.063 0.576 0.081 ;
			RECT 0.234 0.063 0.393 0.081 ;
			RECT 0.234 0.027 0.252 0.081 ;
			RECT 0.146 0.027 0.252 0.045 ;
			RECT 0.308 0.027 0.556 0.045 ;

	END

END OA332x1_ASAP7_75t_L

MACRO OA332x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA332x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.137 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.18 0.225 0.63 0.243 ;
			RECT 0.612 0.063 0.63 0.243 ;
			RECT 0.18 0.189 0.198 0.243 ;
			RECT 0.126 0.189 0.198 0.207 ;
			RECT 0.126 0.119 0.144 0.207 ;
			RECT 0.525 0.063 0.63 0.081 ;
			RECT 0.288 0.063 0.447 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.2 0.027 0.306 0.045 ;
			RECT 0.362 0.027 0.61 0.045 ;

	END

END OA332x2_ASAP7_75t_L

MACRO OA333x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA333x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.63 0.243 ;
			RECT 0.612 0.063 0.63 0.243 ;
			RECT 0.099 0.186 0.117 0.243 ;
			RECT 0.072 0.186 0.117 0.204 ;
			RECT 0.072 0.115 0.09 0.204 ;
			RECT 0.467 0.063 0.63 0.081 ;
			RECT 0.232 0.063 0.394 0.081 ;
			RECT 0.232 0.027 0.25 0.081 ;
			RECT 0.147 0.027 0.25 0.045 ;
			RECT 0.309 0.027 0.569 0.045 ;

	END

END OA333x1_ASAP7_75t_L

MACRO OA333x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA333x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 0.122 0.243 ;
			RECT 0.072 0.027 0.122 0.045 ;
			RECT 0.072 0.027 0.09 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.106 0.63 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.684 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.153 0.186 0.171 0.243 ;
			RECT 0.126 0.186 0.171 0.204 ;
			RECT 0.126 0.115 0.144 0.204 ;
			RECT 0.521 0.063 0.684 0.081 ;
			RECT 0.286 0.063 0.448 0.081 ;
			RECT 0.286 0.027 0.304 0.081 ;
			RECT 0.201 0.027 0.304 0.045 ;
			RECT 0.363 0.027 0.623 0.045 ;

	END

END OA333x2_ASAP7_75t_L

MACRO OA33x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OA33x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.225 0.117 0.243 ;
			RECT 0.099 0.189 0.117 0.243 ;
			RECT 0.062 0.189 0.117 0.207 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.144 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.144 0.126 0.162 0.243 ;
			RECT 0.121 0.126 0.162 0.144 ;
			RECT 0.364 0.063 0.522 0.081 ;
			RECT 0.202 0.027 0.446 0.045 ;

	END

END OA33x2_ASAP7_75t_L

MACRO OAI211xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI211xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.099 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI211xp5_ASAP7_75t_L

MACRO OAI21x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI21x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.369 0.027 0.414 0.045 ;
			RECT 0.018 0.027 0.063 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.189 0.306 0.207 ;
			RECT 0.288 0.106 0.306 0.207 ;
			RECT 0.126 0.106 0.144 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.19 0.127 0.256 0.145 ;
			RECT 0.19 0.099 0.227 0.171 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.072 0.063 0.36 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.027 0.333 0.045 ;

	END

END OAI21x1_ASAP7_75t_L

MACRO OAI21xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI21xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.099 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.203 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI21xp33_ASAP7_75t_L

MACRO OAI21xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI21xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.099 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.203 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI21xp5_ASAP7_75t_L

MACRO OAI221xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI221xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.23 0.243 ;
			RECT 0.018 0.063 0.123 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.201 0.063 0.339 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI221xp5_ASAP7_75t_L

MACRO OAI222xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI222xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.522 0.243 ;
			RECT 0.504 0.055 0.522 0.243 ;
			RECT 0.018 0.063 0.122 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.063 0.36 0.081 ;
			RECT 0.342 0.027 0.36 0.081 ;
			RECT 0.342 0.027 0.468 0.045 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI222xp33_ASAP7_75t_L

MACRO OAI22x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI22x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.038 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.309 0.063 0.522 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.153 0.379 0.171 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.189 0.468 0.207 ;
			RECT 0.45 0.099 0.468 0.207 ;
			RECT 0.431 0.099 0.468 0.117 ;
			RECT 0.288 0.118 0.306 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.161 0.153 0.198 0.171 ;
			RECT 0.18 0.063 0.198 0.171 ;
			RECT 0.161 0.063 0.198 0.081 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.189 0.252 0.207 ;
			RECT 0.234 0.116 0.252 0.207 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.207 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.5 0.045 ;

	END

END OAI22x1_ASAP7_75t_L

MACRO OAI22xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI22xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.063 0.117 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.225 0.275 0.243 ;
			RECT 0.234 0.07 0.252 0.243 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI22xp33_ASAP7_75t_L

MACRO OAI22xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI22xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.063 0.117 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.225 0.275 0.243 ;
			RECT 0.234 0.07 0.252 0.243 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.063 0.198 0.164 ;
			RECT 0.151 0.063 0.198 0.081 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI22xp5_ASAP7_75t_L

MACRO OAI311xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI311xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.198 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END B1
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.027 0.234 0.045 ;

	END

END OAI311xp33_ASAP7_75t_L

MACRO OAI31xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI31xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.256 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.093 0.027 0.23 0.045 ;

	END

END OAI31xp33_ASAP7_75t_L

MACRO OAI31xp67_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI31xp67_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.063 0.663 0.081 ;
			RECT 0.202 0.189 0.252 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.666 0.126 0.684 0.198 ;
			RECT 0.553 0.126 0.684 0.144 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.126 0.419 0.144 ;
			RECT 0.288 0.126 0.306 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.225 0.663 0.243 ;
			RECT 0.364 0.189 0.608 0.207 ;
			RECT 0.04 0.027 0.554 0.045 ;
			RECT 0.094 0.225 0.446 0.243 ;

	END

END OAI31xp67_ASAP7_75t_L

MACRO OAI321xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI321xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.198 0.225 0.414 0.243 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.31 0.063 0.414 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.396 0.045 ;
			RECT 0.094 0.063 0.23 0.081 ;

	END

END OAI321xp33_ASAP7_75t_L

MACRO OAI322xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI322xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.147 0.225 0.468 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.364 0.063 0.468 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.105 0.306 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.105 0.36 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.027 0.45 0.045 ;
			RECT 0.039 0.063 0.284 0.081 ;

	END

END OAI322xp33_ASAP7_75t_L

MACRO OAI32xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI32xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.36 0.243 ;
			RECT 0.342 0.063 0.36 0.243 ;
			RECT 0.256 0.063 0.36 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.063 0.222 0.081 ;
			RECT 0.18 0.063 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.027 0.338 0.045 ;

	END

END OAI32xp33_ASAP7_75t_L

MACRO OAI331xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI331xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.468 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.417 0.063 0.468 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.393 0.045 ;
			RECT 0.092 0.063 0.339 0.081 ;

	END

END OAI331xp33_ASAP7_75t_L

MACRO OAI332xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI332xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.417 0.063 0.522 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.502 0.045 ;
			RECT 0.092 0.063 0.339 0.081 ;

	END

END OAI332xp33_ASAP7_75t_L

MACRO OAI333xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI333xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.413 0.063 0.576 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.515 0.045 ;
			RECT 0.094 0.063 0.34 0.081 ;

	END

END OAI333xp33_ASAP7_75t_L

MACRO OAI33xp33_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OAI33xp33_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.414 0.243 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.256 0.063 0.414 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.092 0.027 0.338 0.045 ;

	END

END OAI33xp33_ASAP7_75t_L

MACRO OR2x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR2x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.207 0.027 0.306 0.045 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.077 0.144 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.186 0.243 ;
			RECT 0.168 0.027 0.186 0.243 ;
			RECT 0.168 0.126 0.227 0.144 ;
			RECT 0.094 0.027 0.186 0.045 ;

	END

END OR2x2_ASAP7_75t_L

MACRO OR2x4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR2x4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.207 0.027 0.414 0.045 ;
			RECT 0.315 0.184 0.333 0.243 ;
			RECT 0.315 0.027 0.333 0.086 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.077 0.144 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.187 0.243 ;
			RECT 0.169 0.027 0.187 0.243 ;
			RECT 0.169 0.126 0.227 0.144 ;
			RECT 0.094 0.027 0.187 0.045 ;

	END

END OR2x4_ASAP7_75t_L

MACRO OR2x6_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR2x6_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.31 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.063 0.144 0.122 ;
			RECT 0.018 0.063 0.144 0.081 ;
			RECT 0.018 0.063 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.153 0.252 0.171 ;
			RECT 0.234 0.121 0.252 0.171 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.189 0.306 0.207 ;
			RECT 0.288 0.07 0.306 0.207 ;
			RECT 0.234 0.07 0.306 0.088 ;
			RECT 0.234 0.027 0.252 0.088 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END OR2x6_ASAP7_75t_L

MACRO OR3x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR3x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.183 0.306 0.201 ;
			RECT 0.288 0.076 0.306 0.201 ;
			RECT 0.261 0.076 0.306 0.094 ;
			RECT 0.261 0.183 0.279 0.235 ;
			RECT 0.261 0.034 0.279 0.094 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.262 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END OR3x1_ASAP7_75t_L

MACRO OR3x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR3x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.261 0.027 0.36 0.045 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.24 0.243 ;
			RECT 0.222 0.027 0.24 0.243 ;
			RECT 0.222 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.24 0.045 ;

	END

END OR3x2_ASAP7_75t_L

MACRO OR3x4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR3x4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.261 0.027 0.468 0.045 ;
			RECT 0.369 0.184 0.387 0.243 ;
			RECT 0.369 0.027 0.387 0.086 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.241 0.243 ;
			RECT 0.223 0.027 0.241 0.243 ;
			RECT 0.223 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.241 0.045 ;

	END

END OR3x4_ASAP7_75t_L

MACRO OR4x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR4x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.072 0.066 0.09 0.152 ;
			RECT 0.072 0.066 0.117 0.084 ;
			RECT 0.099 0.027 0.117 0.084 ;
			RECT 0.099 0.027 0.36 0.045 ;

	END

END OR4x1_ASAP7_75t_L

MACRO OR4x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR4x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.364 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.099 0.063 0.117 0.149 ;
			RECT 0.099 0.063 0.171 0.081 ;
			RECT 0.153 0.027 0.171 0.081 ;
			RECT 0.153 0.027 0.414 0.045 ;

	END

END OR4x2_ASAP7_75t_L

MACRO OR5x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR5x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.35 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.349 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.07 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.288 0.063 0.36 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.018 0.027 0.306 0.045 ;

	END

END OR5x1_ASAP7_75t_L

MACRO OR5x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN OR5x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.343 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.07 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.288 0.063 0.36 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.018 0.027 0.306 0.045 ;

	END

END OR5x2_ASAP7_75t_L

MACRO SDFHx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFHx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.332 0.243 ;
			RECT 1.314 0.027 1.332 0.243 ;
			RECT 1.282 0.027 1.332 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.185 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.185 0.117 0.203 ;
			RECT 0.072 0.081 0.09 0.203 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.284 0.108 0.436 0.126 ;
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.164 ;
			LAYER V1 ;
			RECT 0.396 0.108 0.414 0.126 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.467 0.108 0.59 0.126 ;
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;
			LAYER V1 ;
			RECT 0.504 0.108 0.522 0.126 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.797 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.021 0.225 0.068 0.243 ;
			RECT 0.021 0.027 0.039 0.243 ;
			RECT 0.021 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.016 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.021 0.144 0.039 0.162 ;

	END

END SDFHx1_ASAP7_75t_L

MACRO SDFHx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFHx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.282 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.019 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx2_ASAP7_75t_L

MACRO SDFHx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFHx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.458 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.44 0.243 ;
			RECT 1.422 0.027 1.44 0.243 ;
			RECT 1.282 0.027 1.44 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.458 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.458 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.019 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx3_ASAP7_75t_L

MACRO SDFHx4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFHx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.674 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.444 0.225 1.656 0.243 ;
			RECT 1.637 0.027 1.656 0.243 ;
			RECT 1.444 0.027 1.656 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.164 ;
			RECT 0.378 0.225 0.459 0.243 ;
			RECT 0.378 0.099 0.468 0.117 ;
			RECT 0.378 0.099 0.396 0.243 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.599 0.081 ;
			RECT 0.558 0.063 0.576 0.164 ;
			RECT 0.234 0.126 0.289 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;
			LAYER V1 ;
			RECT 0.234 0.072 0.252 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.027 0.767 0.045 ;
			RECT 0.639 0.063 0.711 0.081 ;
			RECT 0.693 0.027 0.711 0.081 ;
			RECT 0.612 0.106 0.657 0.124 ;
			RECT 0.639 0.063 0.657 0.124 ;
			RECT 0.612 0.106 0.63 0.164 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.674 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.674 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.059 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.368 0.126 1.447 0.144 ;
			RECT 1.242 0.126 1.283 0.144 ;
			RECT 1.242 0.027 1.26 0.144 ;
			RECT 1.113 0.027 1.386 0.045 ;
			RECT 1.206 0.182 1.332 0.2 ;
			RECT 1.314 0.081 1.332 0.2 ;
			RECT 1.206 0.106 1.224 0.2 ;
			RECT 1.287 0.081 1.332 0.099 ;
			RECT 0.882 0.063 0.9 0.164 ;
			RECT 0.882 0.063 0.981 0.081 ;
			RECT 0.801 0.225 0.954 0.243 ;
			RECT 0.936 0.106 0.954 0.243 ;
			RECT 0.801 0.189 0.819 0.243 ;
			RECT 0.738 0.189 0.819 0.207 ;
			RECT 0.738 0.07 0.756 0.207 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.504 0.063 0.522 0.164 ;
			RECT 0.342 0.063 0.522 0.081 ;
			RECT 0.31 0.027 0.36 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.126 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.09 0.045 ;
			RECT 1.152 0.106 1.17 0.2 ;
			RECT 1.098 0.07 1.116 0.164 ;
			RECT 1.044 0.106 1.062 0.2 ;
			RECT 0.828 0.07 0.846 0.167 ;
			RECT 0.774 0.07 0.792 0.164 ;
			RECT 0.58 0.225 0.77 0.243 ;
			RECT 0.684 0.121 0.702 0.167 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.423 0.189 0.662 0.207 ;
			RECT 0.126 0.106 0.144 0.2 ;
			LAYER M2 ;
			RECT 0.019 0.144 1.175 0.162 ;
			RECT 0.175 0.108 1.121 0.126 ;
			LAYER V1 ;
			RECT 1.152 0.144 1.17 0.162 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 1.044 0.144 1.062 0.162 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.108 0.792 0.126 ;
			RECT 0.684 0.144 0.702 0.162 ;
			RECT 0.18 0.108 0.198 0.126 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx4_ASAP7_75t_L

MACRO SDFLx1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFLx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.332 0.243 ;
			RECT 1.314 0.027 1.332 0.243 ;
			RECT 1.282 0.027 1.332 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.797 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx1_ASAP7_75t_L

MACRO SDFLx2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFLx2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.282 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx2_ASAP7_75t_L

MACRO SDFLx3_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFLx3_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.458 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.44 0.243 ;
			RECT 1.422 0.027 1.44 0.243 ;
			RECT 1.282 0.027 1.44 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.458 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.458 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx3_ASAP7_75t_L

MACRO SDFLx4_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN SDFLx4_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.674 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.444 0.225 1.656 0.243 ;
			RECT 1.637 0.027 1.656 0.243 ;
			RECT 1.444 0.027 1.656 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.164 ;
			RECT 0.378 0.225 0.459 0.243 ;
			RECT 0.378 0.099 0.468 0.117 ;
			RECT 0.378 0.099 0.396 0.243 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.599 0.081 ;
			RECT 0.558 0.063 0.576 0.164 ;
			RECT 0.234 0.126 0.289 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;
			LAYER V1 ;
			RECT 0.234 0.072 0.252 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.027 0.767 0.045 ;
			RECT 0.639 0.063 0.711 0.081 ;
			RECT 0.693 0.027 0.711 0.081 ;
			RECT 0.612 0.106 0.657 0.124 ;
			RECT 0.639 0.063 0.657 0.124 ;
			RECT 0.612 0.106 0.63 0.164 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.674 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.674 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.059 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.368 0.126 1.447 0.144 ;
			RECT 1.242 0.126 1.283 0.144 ;
			RECT 1.242 0.027 1.26 0.144 ;
			RECT 1.113 0.027 1.386 0.045 ;
			RECT 1.206 0.182 1.332 0.2 ;
			RECT 1.314 0.081 1.332 0.2 ;
			RECT 1.206 0.106 1.224 0.2 ;
			RECT 1.287 0.081 1.332 0.099 ;
			RECT 0.882 0.063 0.9 0.164 ;
			RECT 0.882 0.063 0.981 0.081 ;
			RECT 0.801 0.225 0.954 0.243 ;
			RECT 0.936 0.106 0.954 0.243 ;
			RECT 0.801 0.189 0.819 0.243 ;
			RECT 0.738 0.189 0.819 0.207 ;
			RECT 0.738 0.07 0.756 0.207 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.504 0.063 0.522 0.164 ;
			RECT 0.342 0.063 0.522 0.081 ;
			RECT 0.31 0.027 0.36 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.126 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.108 0.047 0.126 ;
			RECT 0.009 0.027 0.09 0.045 ;
			RECT 1.152 0.106 1.17 0.2 ;
			RECT 1.098 0.07 1.116 0.164 ;
			RECT 1.044 0.106 1.062 0.2 ;
			RECT 0.828 0.07 0.846 0.167 ;
			RECT 0.774 0.07 0.792 0.164 ;
			RECT 0.58 0.225 0.77 0.243 ;
			RECT 0.684 0.121 0.702 0.167 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.423 0.189 0.662 0.207 ;
			RECT 0.126 0.103 0.144 0.2 ;
			LAYER M2 ;
			RECT 0.175 0.144 1.175 0.162 ;
			RECT 0.019 0.108 1.121 0.126 ;
			LAYER V1 ;
			RECT 1.152 0.144 1.17 0.162 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 1.044 0.144 1.062 0.162 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.108 0.792 0.126 ;
			RECT 0.684 0.144 0.702 0.162 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.108 0.144 0.126 ;
			RECT 0.024 0.108 0.042 0.126 ;

	END

END SDFLx4_ASAP7_75t_L

MACRO TAPCELL_ASAP7_75t_L
	CLASS CORE WELLTAP ;
	FOREIGN TAPCELL_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.108 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.108 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.108 0.279 ;

		END 

	END VDD

END TAPCELL_ASAP7_75t_L

MACRO TAPCELL_WITH_FILLER_ASAP7_75t_L
	CLASS CORE WELLTAP ;
	FOREIGN TAPCELL_WITH_FILLER_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END TAPCELL_WITH_FILLER_ASAP7_75t_L

MACRO TIEHIx1_ASAP7_75t_L
	CLASS CORE TIEHIGH ;
	FOREIGN TIEHIx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN H
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.07 0.144 0.243 ;
			RECT 0.067 0.07 0.144 0.088 ;

		END 

	END H
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.155 0.095 0.173 ;
			RECT 0.018 0.027 0.036 0.173 ;
			RECT 0.018 0.027 0.068 0.045 ;

	END

END TIEHIx1_ASAP7_75t_L

MACRO TIELOx1_ASAP7_75t_L
	CLASS CORE TIELOW ;
	FOREIGN TIELOx1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN L
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.067 0.182 0.144 0.2 ;
			RECT 0.126 0.027 0.144 0.2 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END L
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.097 0.036 0.243 ;
			RECT 0.018 0.097 0.095 0.115 ;

	END

END TIELOx1_ASAP7_75t_L

MACRO XNOR2x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN XNOR2x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.612 0.243 ;
			RECT 0.45 0.077 0.468 0.243 ;
			RECT 0.418 0.077 0.468 0.095 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.121 0.18 0.581 0.198 ;
			LAYER M1 ;
			RECT 0.526 0.189 0.576 0.207 ;
			RECT 0.558 0.121 0.576 0.207 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			LAYER V1 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.558 0.18 0.576 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.298 0.072 0.527 0.09 ;
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.152 ;
			RECT 0.305 0.126 0.365 0.144 ;
			RECT 0.305 0.067 0.323 0.144 ;
			RECT 0.213 0.067 0.323 0.085 ;
			RECT 0.213 0.027 0.231 0.085 ;
			RECT 0.018 0.027 0.231 0.045 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.027 0.036 0.236 ;
			LAYER V1 ;
			RECT 0.305 0.072 0.323 0.09 ;
			RECT 0.504 0.072 0.522 0.09 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.092 0.225 0.193 0.243 ;
			RECT 0.174 0.189 0.193 0.243 ;
			RECT 0.174 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.174 0.082 0.192 0.243 ;
			RECT 0.256 0.027 0.608 0.045 ;

	END

END XNOR2x1_ASAP7_75t_L

MACRO XNOR2x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN XNOR2x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.472 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.44 0.243 ;
			RECT 0.422 0.126 0.44 0.243 ;
			RECT 0.391 0.126 0.44 0.144 ;
			RECT 0.261 0.183 0.279 0.243 ;
			RECT 0.126 0.183 0.279 0.201 ;
			RECT 0.126 0.12 0.144 0.201 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.189 0.38 0.207 ;
			RECT 0.342 0.107 0.36 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.063 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.477 0.063 0.495 0.151 ;
			RECT 0.423 0.063 0.495 0.081 ;
			RECT 0.423 0.027 0.441 0.081 ;
			RECT 0.018 0.027 0.441 0.045 ;
			RECT 0.302 0.063 0.32 0.195 ;
			RECT 0.072 0.063 0.09 0.149 ;
			RECT 0.072 0.063 0.392 0.081 ;
			RECT 0.099 0.225 0.23 0.243 ;

	END

END XNOR2x2_ASAP7_75t_L

MACRO XNOR2xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN XNOR2xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.423 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.207 0.063 0.36 0.081 ;
			RECT 0.207 0.027 0.225 0.081 ;
			RECT 0.072 0.027 0.225 0.045 ;
			RECT 0.072 0.027 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.075 0.18 0.243 ;
			RECT 0.162 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.261 0.027 0.387 0.045 ;

	END

END XNOR2xp5_ASAP7_75t_L

MACRO XOR2x1_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN XOR2x1_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.027 0.612 0.045 ;
			RECT 0.418 0.175 0.468 0.193 ;
			RECT 0.45 0.027 0.468 0.193 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.298 0.18 0.527 0.198 ;
			LAYER M1 ;
			RECT 0.504 0.118 0.522 0.2 ;
			RECT 0.305 0.126 0.365 0.144 ;
			RECT 0.213 0.185 0.323 0.203 ;
			RECT 0.305 0.126 0.323 0.203 ;
			RECT 0.018 0.225 0.231 0.243 ;
			RECT 0.213 0.185 0.231 0.243 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.243 ;
			LAYER V1 ;
			RECT 0.305 0.18 0.323 0.198 ;
			RECT 0.504 0.18 0.522 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.121 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.576 0.149 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.126 0.063 0.144 0.149 ;
			RECT 0.107 0.063 0.144 0.081 ;
			LAYER V1 ;
			RECT 0.126 0.072 0.144 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.174 0.027 0.192 0.188 ;
			RECT 0.396 0.063 0.414 0.149 ;
			RECT 0.174 0.063 0.414 0.081 ;
			RECT 0.174 0.027 0.193 0.081 ;
			RECT 0.092 0.027 0.193 0.045 ;
			RECT 0.256 0.225 0.608 0.243 ;

	END

END XOR2x1_ASAP7_75t_L

MACRO XOR2x2_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN XOR2x2_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.472 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.38 0.081 ;
			RECT 0.342 0.063 0.36 0.163 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.422 0.027 0.44 0.163 ;
			RECT 0.391 0.126 0.44 0.144 ;
			RECT 0.261 0.027 0.44 0.045 ;
			RECT 0.126 0.069 0.279 0.087 ;
			RECT 0.261 0.027 0.279 0.087 ;
			RECT 0.126 0.069 0.144 0.15 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.441 0.243 ;
			RECT 0.423 0.189 0.441 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.423 0.189 0.495 0.207 ;
			RECT 0.477 0.119 0.495 0.207 ;
			RECT 0.018 0.027 0.063 0.045 ;
			RECT 0.072 0.189 0.392 0.207 ;
			RECT 0.302 0.075 0.32 0.207 ;
			RECT 0.072 0.121 0.09 0.207 ;
			RECT 0.099 0.027 0.23 0.045 ;

	END

END XOR2x2_ASAP7_75t_L

MACRO XOR2xp5_ASAP7_75t_L
	CLASS CORE ;
	FOREIGN XOR2xp5_ASAP7_75t_L 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.423 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.256 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.189 0.36 0.207 ;
			RECT 0.342 0.12 0.36 0.207 ;
			RECT 0.018 0.225 0.225 0.243 ;
			RECT 0.207 0.189 0.225 0.243 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.106 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.162 0.027 0.18 0.195 ;
			RECT 0.396 0.063 0.414 0.149 ;
			RECT 0.162 0.063 0.414 0.081 ;
			RECT 0.094 0.027 0.18 0.045 ;
			RECT 0.256 0.225 0.387 0.243 ;

	END

END XOR2xp5_ASAP7_75t_L

MACRO A2O1A1Ixp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN A2O1A1Ixp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.214 0.215 0.306 0.233 ;
			RECT 0.288 0.037 0.306 0.233 ;
			RECT 0.262 0.037 0.306 0.055 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.081 0.252 0.19 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.23 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END A2O1A1Ixp33_ASAP7_75t_SL

MACRO A2O1A1O1Ixp25_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN A2O1A1O1Ixp25_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.423 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.261 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.127 0.414 0.145 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.207 0.225 0.387 0.243 ;
			RECT 0.04 0.027 0.225 0.045 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END A2O1A1O1Ixp25_ASAP7_75t_SL

MACRO AND2x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND2x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.207 0.027 0.306 0.045 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.027 0.18 0.243 ;
			RECT 0.162 0.126 0.203 0.144 ;
			RECT 0.07 0.027 0.088 0.086 ;
			RECT 0.07 0.027 0.18 0.045 ;

	END

END AND2x2_ASAP7_75t_SL

MACRO AND2x4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND2x4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.31 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.028 0.252 0.15 ;
			RECT 0.072 0.028 0.252 0.046 ;
			RECT 0.072 0.028 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.107 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.231 0.243 ;
			RECT 0.18 0.064 0.198 0.243 ;
			RECT 0.179 0.182 0.306 0.2 ;
			RECT 0.288 0.121 0.306 0.2 ;
			RECT 0.115 0.064 0.198 0.082 ;

	END

END AND2x4_ASAP7_75t_SL

MACRO AND2x6_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND2x6_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.554 0.243 ;
			RECT 0.31 0.027 0.554 0.045 ;
			RECT 0.45 0.027 0.468 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.028 0.252 0.15 ;
			RECT 0.072 0.028 0.252 0.046 ;
			RECT 0.072 0.028 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.107 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.231 0.243 ;
			RECT 0.18 0.064 0.198 0.243 ;
			RECT 0.179 0.182 0.306 0.2 ;
			RECT 0.288 0.121 0.306 0.2 ;
			RECT 0.115 0.064 0.198 0.082 ;

	END

END AND2x6_ASAP7_75t_SL

MACRO AND3x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND3x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.183 0.306 0.201 ;
			RECT 0.288 0.076 0.306 0.201 ;
			RECT 0.261 0.076 0.306 0.094 ;
			RECT 0.261 0.183 0.279 0.235 ;
			RECT 0.261 0.034 0.279 0.094 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.263 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END AND3x1_ASAP7_75t_SL

MACRO AND3x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND3x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.261 0.027 0.36 0.045 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END AND3x2_ASAP7_75t_SL

MACRO AND3x4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND3x4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.23 0.243 ;
			RECT 0.018 0.027 0.23 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.189 0.649 0.207 ;
			RECT 0.612 0.099 0.649 0.117 ;
			RECT 0.612 0.099 0.63 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.189 0.541 0.207 ;
			RECT 0.504 0.099 0.541 0.117 ;
			RECT 0.504 0.099 0.522 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.26 0.225 0.746 0.243 ;
			RECT 0.728 0.027 0.746 0.243 ;
			RECT 0.26 0.042 0.278 0.243 ;
			RECT 0.218 0.126 0.278 0.144 ;
			RECT 0.634 0.027 0.746 0.045 ;
			RECT 0.472 0.063 0.701 0.081 ;
			RECT 0.31 0.027 0.554 0.045 ;

	END

END AND3x4_ASAP7_75t_SL

MACRO AND4x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND4x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.299 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.164 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.234 0.189 0.306 0.207 ;
			RECT 0.288 0.12 0.306 0.207 ;
			RECT 0.018 0.027 0.085 0.045 ;

	END

END AND4x1_ASAP7_75t_SL

MACRO AND4x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND4x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.164 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.153 0.189 0.171 0.243 ;
			RECT 0.099 0.189 0.171 0.207 ;
			RECT 0.099 0.119 0.117 0.207 ;
			RECT 0.364 0.027 0.414 0.045 ;

	END

END AND4x2_ASAP7_75t_SL

MACRO AND5x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND5x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.349 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.35 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.164 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.288 0.189 0.36 0.207 ;
			RECT 0.342 0.116 0.36 0.207 ;
			RECT 0.018 0.027 0.07 0.045 ;

	END

END AND5x1_ASAP7_75t_SL

MACRO AND5x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AND5x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.958 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.958 0.027 1.062 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.72 0.189 0.757 0.207 ;
			RECT 0.72 0.099 0.757 0.117 ;
			RECT 0.72 0.099 0.738 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.593 0.189 0.63 0.207 ;
			RECT 0.612 0.099 0.63 0.207 ;
			RECT 0.593 0.099 0.63 0.117 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.189 0.487 0.207 ;
			RECT 0.45 0.099 0.487 0.117 ;
			RECT 0.45 0.099 0.468 0.207 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.269 0.189 0.306 0.207 ;
			RECT 0.288 0.099 0.306 0.207 ;
			RECT 0.269 0.099 0.306 0.117 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.225 0.9 0.243 ;
			RECT 0.882 0.027 0.9 0.243 ;
			RECT 0.882 0.126 0.942 0.144 ;
			RECT 0.742 0.027 0.9 0.045 ;
			RECT 0.58 0.063 0.824 0.081 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.256 0.063 0.5 0.081 ;
			RECT 0.094 0.027 0.338 0.045 ;

	END

END AND5x2_ASAP7_75t_SL

MACRO AO211x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO211x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.742 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.311 0.144 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.215 0.063 0.252 0.081 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.153 0.541 0.171 ;
			RECT 0.504 0.063 0.522 0.171 ;
			RECT 0.485 0.063 0.522 0.081 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.666 0.125 0.743 0.143 ;
			RECT 0.094 0.027 0.684 0.045 ;
			RECT 0.31 0.189 0.608 0.207 ;
			RECT 0.04 0.225 0.393 0.243 ;

	END

END AO211x2_ASAP7_75t_SL

MACRO AO21x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO21x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.23 0.225 0.295 0.243 ;
			RECT 0.277 0.038 0.295 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.189 0.252 0.207 ;
			RECT 0.234 0.027 0.252 0.207 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AO21x1_ASAP7_75t_SL

MACRO AO21x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO21x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.23 0.225 0.333 0.243 ;
			RECT 0.315 0.069 0.333 0.243 ;
			RECT 0.276 0.069 0.333 0.087 ;
			RECT 0.276 0.038 0.294 0.087 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.189 0.252 0.207 ;
			RECT 0.234 0.027 0.252 0.207 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AO21x2_ASAP7_75t_SL

MACRO AO221x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO221x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.459 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.126 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;
			RECT 0.396 0.126 0.474 0.144 ;
			RECT 0.396 0.027 0.414 0.144 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.2 0.189 0.339 0.207 ;
			RECT 0.039 0.225 0.176 0.243 ;

	END

END AO221x1_ASAP7_75t_SL

MACRO AO221x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO221x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.549 0.243 ;
			RECT 0.531 0.027 0.549 0.243 ;
			RECT 0.459 0.027 0.549 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.126 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;
			RECT 0.396 0.126 0.474 0.144 ;
			RECT 0.396 0.027 0.414 0.144 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.2 0.189 0.339 0.207 ;
			RECT 0.039 0.225 0.176 0.243 ;

	END

END AO221x2_ASAP7_75t_SL

MACRO AO222x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO222x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.526 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.531 0.027 0.63 0.045 ;
			RECT 0.531 0.027 0.549 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.009 0.189 0.122 0.207 ;
			RECT 0.009 0.027 0.027 0.207 ;
			RECT 0.486 0.126 0.554 0.144 ;
			RECT 0.486 0.027 0.504 0.144 ;
			RECT 0.009 0.027 0.504 0.045 ;
			RECT 0.342 0.225 0.468 0.243 ;
			RECT 0.342 0.189 0.36 0.243 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO222x2_ASAP7_75t_SL

MACRO AO22x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO22x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.418 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.287 0.081 ;
			RECT 0.234 0.063 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.342 0.126 0.419 0.144 ;
			RECT 0.107 0.027 0.36 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO22x1_ASAP7_75t_SL

MACRO AO22x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO22x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.418 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.287 0.081 ;
			RECT 0.234 0.063 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.342 0.126 0.419 0.144 ;
			RECT 0.107 0.027 0.36 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AO22x2_ASAP7_75t_SL

MACRO AO31x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO31x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.741 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.742 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.099 0.576 0.149 ;
			RECT 0.504 0.099 0.576 0.117 ;
			RECT 0.485 0.153 0.522 0.171 ;
			RECT 0.504 0.099 0.522 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.414 0.149 ;
			RECT 0.288 0.099 0.414 0.117 ;
			RECT 0.288 0.153 0.325 0.171 ;
			RECT 0.288 0.07 0.306 0.171 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.059 0.207 ;
			RECT 0.018 0.027 0.059 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.612 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.612 0.189 0.63 0.243 ;
			RECT 0.199 0.189 0.63 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.666 0.126 0.797 0.144 ;
			RECT 0.2 0.063 0.252 0.081 ;
			RECT 0.526 0.027 0.684 0.045 ;
			RECT 0.364 0.063 0.608 0.081 ;
			RECT 0.04 0.225 0.554 0.243 ;
			RECT 0.094 0.027 0.447 0.045 ;

	END

END AO31x2_ASAP7_75t_SL

MACRO AO322x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO322x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.634 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.634 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.153 0.325 0.171 ;
			RECT 0.288 0.063 0.325 0.081 ;
			RECT 0.288 0.063 0.306 0.171 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.063 0.541 0.081 ;
			RECT 0.504 0.063 0.522 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.396 0.189 0.576 0.207 ;
			RECT 0.558 0.126 0.576 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.558 0.126 0.743 0.144 ;
			RECT 0.04 0.027 0.446 0.045 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.189 0.198 0.243 ;
			RECT 0.18 0.189 0.338 0.207 ;
			RECT 0.256 0.225 0.5 0.243 ;

	END

END AO322x2_ASAP7_75t_SL

MACRO AO32x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO32x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.063 0.063 0.081 ;
			RECT 0.045 0.034 0.063 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.062 0.126 0.108 0.144 ;
			RECT 0.09 0.027 0.108 0.144 ;
			RECT 0.09 0.027 0.414 0.045 ;
			RECT 0.148 0.225 0.392 0.243 ;

	END

END AO32x1_ASAP7_75t_SL

MACRO AO32x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO32x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.068 0.117 0.086 ;
			RECT 0.099 0.037 0.117 0.086 ;
			RECT 0.018 0.068 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.189 0.33 0.207 ;
			RECT 0.288 0.07 0.306 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.364 0.189 0.468 0.207 ;
			RECT 0.45 0.027 0.468 0.207 ;
			RECT 0.093 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.468 0.045 ;
			RECT 0.202 0.225 0.446 0.243 ;

	END

END AO32x2_ASAP7_75t_SL

MACRO AO331x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO331x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.081 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B3
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.072 0.063 0.09 0.152 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.522 0.045 ;
			RECT 0.308 0.189 0.447 0.207 ;
			RECT 0.146 0.225 0.393 0.243 ;

	END

END AO331x1_ASAP7_75t_SL

MACRO AO331x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO331x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.027 0.135 0.045 ;
			RECT 0.072 0.225 0.122 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.126 0.063 0.144 0.152 ;
			RECT 0.126 0.063 0.198 0.081 ;
			RECT 0.18 0.027 0.198 0.081 ;
			RECT 0.18 0.027 0.576 0.045 ;
			RECT 0.362 0.189 0.501 0.207 ;
			RECT 0.2 0.225 0.447 0.243 ;

	END

END AO331x2_ASAP7_75t_SL

MACRO AO332x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO332x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.094 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.072 0.063 0.09 0.151 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.576 0.045 ;
			RECT 0.146 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.234 0.189 0.393 0.207 ;
			RECT 0.308 0.225 0.556 0.243 ;

	END

END AO332x1_ASAP7_75t_SL

MACRO AO332x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO332x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.148 0.045 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.189 0.63 0.207 ;
			RECT 0.612 0.027 0.63 0.207 ;
			RECT 0.126 0.063 0.144 0.151 ;
			RECT 0.126 0.063 0.198 0.081 ;
			RECT 0.18 0.027 0.198 0.081 ;
			RECT 0.18 0.027 0.63 0.045 ;
			RECT 0.2 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.288 0.189 0.447 0.207 ;
			RECT 0.362 0.225 0.61 0.243 ;

	END

END AO332x2_ASAP7_75t_SL

MACRO AO333x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO333x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.081 0.045 ;
			RECT 0.018 0.225 0.069 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.471 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.063 0.09 0.152 ;
			RECT 0.072 0.063 0.144 0.081 ;
			RECT 0.126 0.027 0.144 0.081 ;
			RECT 0.126 0.027 0.63 0.045 ;
			RECT 0.31 0.189 0.576 0.207 ;
			RECT 0.148 0.225 0.395 0.243 ;

	END

END AO333x1_ASAP7_75t_SL

MACRO AO333x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO333x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.081 0.117 0.099 ;
			RECT 0.099 0.045 0.117 0.099 ;
			RECT 0.018 0.081 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.07 0.63 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.07 0.576 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.525 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.067 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.684 0.045 ;
			RECT 0.364 0.189 0.63 0.207 ;
			RECT 0.202 0.225 0.449 0.243 ;

	END

END AO333x2_ASAP7_75t_SL

MACRO AO33x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AO33x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.068 0.117 0.086 ;
			RECT 0.099 0.037 0.117 0.086 ;
			RECT 0.018 0.068 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.361 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.067 0.126 0.162 0.144 ;
			RECT 0.144 0.027 0.162 0.144 ;
			RECT 0.144 0.027 0.522 0.045 ;
			RECT 0.199 0.225 0.449 0.243 ;

	END

END AO33x2_ASAP7_75t_SL

MACRO AOI211x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI211x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.519 0.189 0.63 0.207 ;
			RECT 0.612 0.027 0.63 0.207 ;
			RECT 0.091 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.126 0.229 0.144 ;
			RECT 0.18 0.189 0.223 0.207 ;
			RECT 0.18 0.063 0.22 0.081 ;
			RECT 0.18 0.063 0.198 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.123 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.153 0.442 0.171 ;
			RECT 0.396 0.063 0.442 0.081 ;
			RECT 0.396 0.063 0.414 0.171 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.126 0.554 0.144 ;
			RECT 0.504 0.063 0.55 0.081 ;
			RECT 0.504 0.063 0.522 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.306 0.243 ;
			RECT 0.288 0.189 0.306 0.243 ;
			RECT 0.288 0.189 0.449 0.207 ;
			RECT 0.361 0.225 0.608 0.243 ;

	END

END AOI211x1_ASAP7_75t_SL

MACRO AOI211xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI211xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.04 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AOI211xp5_ASAP7_75t_SL

MACRO AOI21x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI21x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.369 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.018 0.027 0.414 0.045 ;
			RECT 0.018 0.225 0.063 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.063 0.306 0.164 ;
			RECT 0.126 0.063 0.306 0.081 ;
			RECT 0.126 0.063 0.144 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.19 0.125 0.256 0.143 ;
			RECT 0.19 0.099 0.227 0.171 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.189 0.36 0.207 ;
			RECT 0.342 0.116 0.36 0.207 ;
			RECT 0.072 0.07 0.09 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.333 0.243 ;

	END

END AOI21x1_ASAP7_75t_SL

MACRO AOI21xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI21xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.107 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END AOI21xp33_ASAP7_75t_SL

MACRO AOI21xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI21xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.142 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.034 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.171 0.243 ;

	END

END AOI21xp5_ASAP7_75t_SL

MACRO AOI221x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI221x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.634 0.189 0.738 0.207 ;
			RECT 0.72 0.045 0.738 0.207 ;
			RECT 0.256 0.045 0.738 0.063 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.153 0.217 0.171 ;
			RECT 0.18 0.027 0.198 0.171 ;
			RECT 0.161 0.027 0.198 0.045 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.126 0.149 0.144 ;
			RECT 0.053 0.153 0.09 0.171 ;
			RECT 0.072 0.027 0.09 0.171 ;
			RECT 0.053 0.027 0.09 0.045 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.081 0.325 0.099 ;
			RECT 0.269 0.153 0.306 0.171 ;
			RECT 0.288 0.081 0.306 0.171 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.153 0.487 0.171 ;
			RECT 0.45 0.081 0.468 0.171 ;
			RECT 0.391 0.126 0.468 0.144 ;
			RECT 0.431 0.081 0.468 0.099 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.126 0.636 0.144 ;
			RECT 0.539 0.189 0.576 0.207 ;
			RECT 0.558 0.081 0.576 0.207 ;
			RECT 0.539 0.081 0.576 0.099 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.225 0.716 0.243 ;
			RECT 0.04 0.189 0.5 0.207 ;

	END

END AOI221x1_ASAP7_75t_SL

MACRO AOI221xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI221xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.23 0.045 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.201 0.189 0.339 0.207 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END AOI221xp5_ASAP7_75t_SL

MACRO AOI222xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI222xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.399 0.045 ;
			RECT 0.018 0.189 0.122 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.034 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.342 0.225 0.468 0.243 ;
			RECT 0.342 0.189 0.36 0.243 ;
			RECT 0.202 0.189 0.36 0.207 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI222xp33_ASAP7_75t_SL

MACRO AOI22x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI22x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.309 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.038 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.153 0.379 0.171 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.431 0.153 0.468 0.171 ;
			RECT 0.45 0.063 0.468 0.171 ;
			RECT 0.288 0.063 0.468 0.081 ;
			RECT 0.288 0.063 0.306 0.152 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.161 0.189 0.198 0.207 ;
			RECT 0.18 0.099 0.198 0.207 ;
			RECT 0.161 0.099 0.198 0.117 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.252 0.154 ;
			RECT 0.072 0.063 0.252 0.081 ;
			RECT 0.072 0.189 0.109 0.207 ;
			RECT 0.072 0.063 0.09 0.207 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.5 0.243 ;

	END

END AOI22x1_ASAP7_75t_SL

MACRO AOI22xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI22xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI22xp33_ASAP7_75t_SL

MACRO AOI22xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI22xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.07 0.144 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END AOI22xp5_ASAP7_75t_SL

MACRO AOI311xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI311xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.198 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.234 0.243 ;

	END

END AOI311xp33_ASAP7_75t_SL

MACRO AOI31xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI31xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.201 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.093 0.225 0.23 0.243 ;

	END

END AOI31xp33_ASAP7_75t_SL

MACRO AOI31xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI31xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.585 0.225 0.663 0.243 ;
			RECT 0.585 0.189 0.603 0.243 ;
			RECT 0.202 0.189 0.603 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;
			RECT 0.202 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.666 0.07 0.684 0.2 ;
			RECT 0.553 0.126 0.684 0.144 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.126 0.419 0.144 ;
			RECT 0.288 0.063 0.325 0.081 ;
			RECT 0.288 0.063 0.306 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.059 0.207 ;
			RECT 0.018 0.027 0.059 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.027 0.663 0.045 ;
			RECT 0.364 0.081 0.608 0.099 ;
			RECT 0.04 0.225 0.554 0.243 ;
			RECT 0.094 0.027 0.447 0.045 ;

	END

END AOI31xp67_ASAP7_75t_SL

MACRO AOI321xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI321xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.198 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.225 0.396 0.243 ;
			RECT 0.094 0.189 0.23 0.207 ;

	END

END AOI321xp33_ASAP7_75t_SL

MACRO AOI322xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI322xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.189 0.468 0.207 ;
			RECT 0.45 0.027 0.468 0.207 ;
			RECT 0.147 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.165 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.165 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.225 0.45 0.243 ;
			RECT 0.039 0.189 0.284 0.207 ;

	END

END AOI322xp5_ASAP7_75t_SL

MACRO AOI32xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI32xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.36 0.207 ;
			RECT 0.342 0.027 0.36 0.207 ;
			RECT 0.04 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.058 0.243 ;
			RECT 0.018 0.063 0.058 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.104 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.104 0.063 0.144 0.081 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.222 0.207 ;
			RECT 0.18 0.07 0.198 0.207 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END AOI32xp33_ASAP7_75t_SL

MACRO AOI331xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI331xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.417 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.201 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.189 0.393 0.207 ;
			RECT 0.092 0.225 0.339 0.243 ;

	END

END AOI331xp33_ASAP7_75t_SL

MACRO AOI332xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI332xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.417 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.201 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.225 0.502 0.243 ;
			RECT 0.092 0.189 0.339 0.207 ;

	END

END AOI332xp33_ASAP7_75t_SL

MACRO AOI333xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI333xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.413 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.201 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.164 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.164 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.164 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.225 0.515 0.243 ;
			RECT 0.094 0.189 0.34 0.207 ;

	END

END AOI333xp33_ASAP7_75t_SL

MACRO AOI33xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN AOI33xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.189 0.414 0.207 ;
			RECT 0.396 0.027 0.414 0.207 ;
			RECT 0.201 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.164 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.338 0.243 ;

	END

END AOI33xp33_ASAP7_75t_SL

MACRO BUFx10_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx10_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.199 0.027 0.738 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.689 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx10_ASAP7_75t_SL

MACRO BUFx12_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx12_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.846 0.243 ;
			RECT 0.828 0.027 0.846 0.243 ;
			RECT 0.199 0.027 0.846 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.8 0.144 ;
			RECT 0.094 0.027 0.144 0.045 ;

	END

END BUFx12_ASAP7_75t_SL

MACRO BUFx12f_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx12f_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.972 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.31 0.027 0.954 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.074 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.972 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.972 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.243 ;
			RECT 0.261 0.126 0.311 0.144 ;
			RECT 0.094 0.027 0.279 0.045 ;

	END

END BUFx12f_ASAP7_75t_SL

MACRO BUFx16f_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx16f_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 1.17 0.243 ;
			RECT 1.152 0.027 1.17 0.243 ;
			RECT 0.31 0.027 1.17 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.06 0.243 ;
			RECT 0.018 0.027 0.06 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.234 0.126 1.124 0.144 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END BUFx16f_ASAP7_75t_SL

MACRO BUFx24_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx24_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.62 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 1.602 0.243 ;
			RECT 1.584 0.027 1.602 0.243 ;
			RECT 0.31 0.027 1.602 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.62 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.62 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.234 0.126 1.553 0.144 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END BUFx24_ASAP7_75t_SL

MACRO BUFx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.145 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.203 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx2_ASAP7_75t_SL

MACRO BUFx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.145 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.26 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx3_ASAP7_75t_SL

MACRO BUFx4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.357 0.243 ;
			RECT 0.339 0.027 0.357 0.243 ;
			RECT 0.145 0.027 0.357 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.314 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx4_ASAP7_75t_SL

MACRO BUFx4f_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx4f_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.199 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.199 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.098 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.367 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx4f_ASAP7_75t_SL

MACRO BUFx5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.145 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.145 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.073 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.12 0.243 ;
			RECT 0.102 0.027 0.12 0.243 ;
			RECT 0.102 0.126 0.368 0.144 ;
			RECT 0.04 0.027 0.12 0.045 ;

	END

END BUFx5_ASAP7_75t_SL

MACRO BUFx6f_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx6f_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.202 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.473 0.144 ;
			RECT 0.094 0.027 0.144 0.045 ;

	END

END BUFx6f_ASAP7_75t_SL

MACRO BUFx8_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN BUFx8_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.202 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.098 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.091 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.581 0.144 ;
			RECT 0.091 0.027 0.144 0.045 ;

	END

END BUFx8_ASAP7_75t_SL

MACRO CKINVDCx10_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx10_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.296 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.224 0.243 ;
			RECT 1.206 0.063 1.224 0.243 ;
			RECT 1.174 0.063 1.224 0.081 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.17 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.296 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.296 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx10_ASAP7_75t_SL

MACRO CKINVDCx11_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx11_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.31 0.243 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.354 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx11_ASAP7_75t_SL

MACRO CKINVDCx12_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx12_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.31 0.243 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.354 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx12_ASAP7_75t_SL

MACRO CKINVDCx14_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx14_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.512 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.44 0.243 ;
			RECT 1.422 0.063 1.44 0.243 ;
			RECT 1.39 0.063 1.44 0.081 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.397 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.512 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.512 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx14_ASAP7_75t_SL

MACRO CKINVDCx16_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx16_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.62 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 1.548 0.243 ;
			RECT 1.53 0.063 1.548 0.243 ;
			RECT 1.498 0.063 1.548 0.081 ;
			RECT 1.368 0.063 1.418 0.081 ;
			RECT 1.368 0.063 1.386 0.243 ;
			RECT 1.098 0.063 1.116 0.243 ;
			RECT 1.066 0.063 1.116 0.081 ;
			RECT 0.936 0.063 0.986 0.081 ;
			RECT 0.936 0.063 0.954 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.634 0.063 0.684 0.081 ;
			RECT 0.504 0.063 0.554 0.081 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.202 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.122 0.081 ;
			RECT 0.072 0.063 0.09 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.412 0.126 1.505 0.144 ;
			RECT 1.444 0.027 1.462 0.144 ;
			RECT 0.158 0.027 1.462 0.045 ;
			RECT 0.98 0.126 1.072 0.144 ;
			RECT 1.017 0.027 1.035 0.144 ;
			RECT 0.547 0.126 0.639 0.144 ;
			RECT 0.584 0.027 0.602 0.144 ;
			RECT 0.126 0.126 0.208 0.144 ;
			RECT 0.158 0.027 0.176 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.62 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.62 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.26 0.126 1.316 0.144 ;
			RECT 1.26 0.09 1.278 0.144 ;
			RECT 1.174 0.09 1.326 0.108 ;
			RECT 1.155 0.162 1.31 0.18 ;
			RECT 1.206 0.126 1.224 0.18 ;
			RECT 1.166 0.126 1.224 0.144 ;
			RECT 0.742 0.162 0.897 0.18 ;
			RECT 0.828 0.126 0.846 0.18 ;
			RECT 0.828 0.126 0.886 0.144 ;
			RECT 0.736 0.126 0.792 0.144 ;
			RECT 0.774 0.09 0.792 0.144 ;
			RECT 0.726 0.09 0.878 0.108 ;
			RECT 0.31 0.162 0.465 0.18 ;
			RECT 0.396 0.126 0.414 0.18 ;
			RECT 0.396 0.126 0.454 0.144 ;
			RECT 0.304 0.126 0.36 0.144 ;
			RECT 0.342 0.09 0.36 0.144 ;
			RECT 0.294 0.09 0.446 0.108 ;

	END

END CKINVDCx16_ASAP7_75t_SL

MACRO CKINVDCx20_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx20_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.052 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 1.98 0.243 ;
			RECT 1.962 0.063 1.98 0.243 ;
			RECT 1.93 0.063 1.98 0.081 ;
			RECT 1.8 0.063 1.85 0.081 ;
			RECT 1.8 0.063 1.818 0.243 ;
			RECT 1.53 0.063 1.548 0.243 ;
			RECT 1.498 0.063 1.548 0.081 ;
			RECT 1.368 0.063 1.418 0.081 ;
			RECT 1.368 0.063 1.386 0.243 ;
			RECT 1.098 0.063 1.116 0.243 ;
			RECT 1.066 0.063 1.116 0.081 ;
			RECT 0.936 0.063 0.986 0.081 ;
			RECT 0.936 0.063 0.954 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.634 0.063 0.684 0.081 ;
			RECT 0.504 0.063 0.554 0.081 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.202 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.122 0.081 ;
			RECT 0.072 0.063 0.09 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.844 0.126 1.937 0.144 ;
			RECT 1.876 0.027 1.894 0.144 ;
			RECT 0.158 0.027 1.894 0.045 ;
			RECT 1.412 0.126 1.505 0.144 ;
			RECT 1.444 0.027 1.462 0.144 ;
			RECT 0.98 0.126 1.072 0.144 ;
			RECT 1.017 0.027 1.035 0.144 ;
			RECT 0.547 0.126 0.639 0.144 ;
			RECT 0.584 0.027 0.602 0.144 ;
			RECT 0.126 0.126 0.208 0.144 ;
			RECT 0.158 0.027 0.176 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.052 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.052 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.692 0.126 1.748 0.144 ;
			RECT 1.692 0.09 1.71 0.144 ;
			RECT 1.606 0.09 1.758 0.108 ;
			RECT 1.587 0.162 1.742 0.18 ;
			RECT 1.638 0.126 1.656 0.18 ;
			RECT 1.598 0.126 1.656 0.144 ;
			RECT 1.26 0.126 1.316 0.144 ;
			RECT 1.26 0.09 1.278 0.144 ;
			RECT 1.174 0.09 1.326 0.108 ;
			RECT 1.155 0.162 1.31 0.18 ;
			RECT 1.206 0.126 1.224 0.18 ;
			RECT 1.166 0.126 1.224 0.144 ;
			RECT 0.742 0.162 0.897 0.18 ;
			RECT 0.828 0.126 0.846 0.18 ;
			RECT 0.828 0.126 0.886 0.144 ;
			RECT 0.736 0.126 0.792 0.144 ;
			RECT 0.774 0.09 0.792 0.144 ;
			RECT 0.726 0.09 0.878 0.108 ;
			RECT 0.31 0.162 0.465 0.18 ;
			RECT 0.396 0.126 0.414 0.18 ;
			RECT 0.396 0.126 0.454 0.144 ;
			RECT 0.304 0.126 0.36 0.144 ;
			RECT 0.342 0.09 0.36 0.144 ;
			RECT 0.294 0.09 0.446 0.108 ;

	END

END CKINVDCx20_ASAP7_75t_SL

MACRO CKINVDCx5p33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx5p33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.094 0.243 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.138 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx5p33_ASAP7_75t_SL

MACRO CKINVDCx6p67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx6p67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.296 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.224 0.243 ;
			RECT 1.206 0.063 1.224 0.243 ;
			RECT 1.174 0.063 1.224 0.081 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.17 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.296 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.296 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx6p67_ASAP7_75t_SL

MACRO CKINVDCx8_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx8_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.094 0.243 ;
			RECT 1.044 0.063 1.094 0.081 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.72 0.063 0.77 0.081 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.418 0.063 0.468 0.081 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.088 0.126 1.138 0.144 ;
			RECT 1.12 0.027 1.138 0.144 ;
			RECT 0.05 0.027 1.138 0.045 ;
			RECT 0.764 0.126 0.814 0.144 ;
			RECT 0.796 0.027 0.814 0.144 ;
			RECT 0.374 0.126 0.424 0.144 ;
			RECT 0.374 0.027 0.392 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.936 0.126 0.992 0.144 ;
			RECT 0.936 0.09 0.954 0.144 ;
			RECT 0.85 0.09 1.002 0.108 ;
			RECT 0.831 0.162 0.986 0.18 ;
			RECT 0.882 0.126 0.9 0.18 ;
			RECT 0.842 0.126 0.9 0.144 ;
			RECT 0.526 0.162 0.681 0.18 ;
			RECT 0.612 0.126 0.63 0.18 ;
			RECT 0.612 0.126 0.67 0.144 ;
			RECT 0.52 0.126 0.576 0.144 ;
			RECT 0.558 0.09 0.576 0.144 ;
			RECT 0.51 0.09 0.662 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx8_ASAP7_75t_SL

MACRO CKINVDCx9p33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN CKINVDCx9p33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.512 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 1.44 0.243 ;
			RECT 1.422 0.063 1.44 0.243 ;
			RECT 1.39 0.063 1.44 0.081 ;
			RECT 1.26 0.063 1.31 0.081 ;
			RECT 1.26 0.063 1.278 0.243 ;
			RECT 0.99 0.063 1.008 0.243 ;
			RECT 0.958 0.063 1.008 0.081 ;
			RECT 0.828 0.063 0.878 0.081 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.396 0.063 0.446 0.081 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.126 0.063 0.144 0.243 ;
			RECT 0.094 0.063 0.144 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 1.304 0.126 1.397 0.144 ;
			RECT 1.336 0.027 1.354 0.144 ;
			RECT 0.05 0.027 1.354 0.045 ;
			RECT 0.872 0.126 0.964 0.144 ;
			RECT 0.909 0.027 0.927 0.144 ;
			RECT 0.439 0.126 0.531 0.144 ;
			RECT 0.476 0.027 0.494 0.144 ;
			RECT 0.05 0.126 0.1 0.144 ;
			RECT 0.05 0.027 0.068 0.144 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.512 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.512 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.126 1.208 0.144 ;
			RECT 1.152 0.09 1.17 0.144 ;
			RECT 1.066 0.09 1.218 0.108 ;
			RECT 1.047 0.162 1.202 0.18 ;
			RECT 1.098 0.126 1.116 0.18 ;
			RECT 1.058 0.126 1.116 0.144 ;
			RECT 0.634 0.162 0.789 0.18 ;
			RECT 0.72 0.126 0.738 0.18 ;
			RECT 0.72 0.126 0.778 0.144 ;
			RECT 0.628 0.126 0.684 0.144 ;
			RECT 0.666 0.09 0.684 0.144 ;
			RECT 0.618 0.09 0.77 0.108 ;
			RECT 0.202 0.162 0.357 0.18 ;
			RECT 0.288 0.126 0.306 0.18 ;
			RECT 0.288 0.126 0.346 0.144 ;
			RECT 0.196 0.126 0.252 0.144 ;
			RECT 0.234 0.09 0.252 0.144 ;
			RECT 0.186 0.09 0.338 0.108 ;

	END

END CKINVDCx9p33_ASAP7_75t_SL

MACRO DECAPx10_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN DECAPx10_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.558 0.045 0.576 0.15 ;
			RECT 0.558 0.045 1.148 0.063 ;
			RECT 0.04 0.207 0.63 0.225 ;
			RECT 0.612 0.121 0.63 0.225 ;

	END

END DECAPx10_ASAP7_75t_SL

MACRO DECAPx1_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN DECAPx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.207 0.144 0.225 ;
			RECT 0.126 0.121 0.144 0.225 ;
			RECT 0.072 0.045 0.09 0.15 ;
			RECT 0.072 0.045 0.122 0.063 ;

	END

END DECAPx1_ASAP7_75t_SL

MACRO DECAPx2_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN DECAPx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.045 0.144 0.15 ;
			RECT 0.126 0.045 0.284 0.063 ;
			RECT 0.04 0.207 0.198 0.225 ;
			RECT 0.18 0.121 0.198 0.225 ;

	END

END DECAPx2_ASAP7_75t_SL

MACRO DECAPx2b_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN DECAPx2b_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.162 0.249 0.18 ;
			RECT 0.18 0.126 0.198 0.18 ;
			RECT 0.18 0.126 0.238 0.144 ;
			RECT 0.088 0.126 0.144 0.144 ;
			RECT 0.126 0.09 0.144 0.144 ;
			RECT 0.078 0.09 0.23 0.108 ;

	END

END DECAPx2b_ASAP7_75t_SL

MACRO DECAPx4_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN DECAPx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.234 0.045 0.252 0.15 ;
			RECT 0.234 0.045 0.5 0.063 ;
			RECT 0.04 0.207 0.306 0.225 ;
			RECT 0.288 0.121 0.306 0.225 ;

	END

END DECAPx4_ASAP7_75t_SL

MACRO DECAPx6_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN DECAPx6_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.342 0.045 0.36 0.15 ;
			RECT 0.342 0.045 0.716 0.063 ;
			RECT 0.04 0.207 0.414 0.225 ;
			RECT 0.396 0.121 0.414 0.225 ;

	END

END DECAPx6_ASAP7_75t_SL

MACRO DFFASRHQNx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFASRHQNx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.336 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.336 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.182 0.117 0.236 ;
			RECT 0.072 0.182 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN RESETN
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.632 0.144 1.067 0.162 ;
			LAYER M1 ;
			RECT 1.044 0.102 1.062 0.167 ;
			RECT 0.612 0.072 0.668 0.09 ;
			RECT 0.612 0.144 0.662 0.162 ;
			RECT 0.612 0.072 0.63 0.162 ;
			LAYER V1 ;
			RECT 0.637 0.144 0.655 0.162 ;
			RECT 1.044 0.144 1.062 0.162 ;

		END 

	END RESETN
	PIN SETN
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.783 0.18 1.067 0.198 ;
			LAYER M1 ;
			RECT 0.774 0.18 0.811 0.198 ;
			RECT 0.774 0.097 0.792 0.198 ;
			LAYER V1 ;
			RECT 0.788 0.18 0.806 0.198 ;

		END 

	END SETN
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.963 0.036 0.981 0.234 ;
			RECT 0.963 0.036 1.008 0.054 ;
			RECT 0.855 0.222 0.936 0.24 ;
			RECT 0.918 0.053 0.936 0.24 ;
			RECT 0.693 0.036 0.711 0.212 ;
			RECT 0.558 0.036 0.576 0.106 ;
			RECT 0.558 0.036 0.77 0.054 ;
			RECT 0.486 0.18 0.547 0.198 ;
			RECT 0.486 0.027 0.504 0.198 ;
			RECT 0.418 0.027 0.504 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.142 0.027 0.198 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.018 0.108 0.047 0.126 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 1.314 0.103 1.332 0.18 ;
			RECT 1.17 0.216 1.202 0.234 ;
			RECT 1.098 0.102 1.116 0.167 ;
			RECT 0.882 0.067 0.9 0.173 ;
			RECT 0.829 0.103 0.847 0.171 ;
			RECT 0.778 0.216 0.819 0.234 ;
			RECT 0.729 0.137 0.747 0.203 ;
			RECT 0.415 0.225 0.608 0.243 ;
			RECT 0.45 0.103 0.468 0.151 ;
			RECT 0.396 0.067 0.414 0.15 ;
			RECT 0.369 0.169 0.387 0.216 ;
			RECT 0.342 0.103 0.36 0.15 ;
			RECT 0.142 0.07 0.16 0.164 ;
			LAYER M2 ;
			RECT 0.913 0.108 1.337 0.126 ;
			RECT 0.783 0.216 1.198 0.234 ;
			RECT 0.741 0.036 1.008 0.054 ;
			RECT 0.018 0.072 0.926 0.09 ;
			RECT 0.175 0.108 0.852 0.126 ;
			RECT 0.364 0.18 0.752 0.198 ;
			LAYER V1 ;
			RECT 1.314 0.108 1.332 0.126 ;
			RECT 1.175 0.216 1.193 0.234 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 0.985 0.036 1.003 0.054 ;
			RECT 0.918 0.108 0.936 0.126 ;
			RECT 0.882 0.072 0.9 0.09 ;
			RECT 0.829 0.108 0.847 0.126 ;
			RECT 0.788 0.216 0.806 0.234 ;
			RECT 0.746 0.036 0.764 0.054 ;
			RECT 0.729 0.18 0.747 0.198 ;
			RECT 0.512 0.18 0.53 0.198 ;
			RECT 0.45 0.108 0.468 0.126 ;
			RECT 0.396 0.072 0.414 0.09 ;
			RECT 0.369 0.18 0.387 0.198 ;
			RECT 0.342 0.108 0.36 0.126 ;
			RECT 0.18 0.108 0.198 0.126 ;
			RECT 0.142 0.072 0.16 0.09 ;
			RECT 0.018 0.072 0.036 0.09 ;

	END

END DFFASRHQNx1_ASAP7_75t_SL

MACRO DFFHQNx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFHQNx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 1.012 0.027 1.062 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx1_ASAP7_75t_SL

MACRO DFFHQNx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFHQNx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.216 1.117 0.234 ;
			RECT 1.099 0.036 1.117 0.234 ;
			RECT 1.012 0.036 1.117 0.054 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx2_ASAP7_75t_SL

MACRO DFFHQNx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFHQNx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.171 0.243 ;
			RECT 1.153 0.027 1.171 0.243 ;
			RECT 1.012 0.027 1.171 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.576 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQNx3_ASAP7_75t_SL

MACRO DFFHQx4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFHQx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.125 0.225 1.333 0.243 ;
			RECT 1.313 0.027 1.333 0.243 ;
			RECT 1.125 0.027 1.333 0.045 ;
			RECT 1.125 0.201 1.143 0.243 ;
			RECT 1.125 0.027 1.143 0.069 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.126 0.29 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.012 0.225 1.098 0.243 ;
			RECT 1.08 0.027 1.098 0.243 ;
			RECT 1.08 0.127 1.175 0.145 ;
			RECT 1.012 0.027 1.098 0.045 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.224 0.738 0.242 ;
			RECT 0.72 0.027 0.738 0.242 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.045 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.315 0.126 0.333 0.203 ;
			RECT 0.315 0.126 0.367 0.144 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.101 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.142 0.106 0.16 0.167 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.019 0.144 0.689 0.162 ;
			RECT 0.175 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.315 0.18 0.333 0.198 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.142 0.144 0.16 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DFFHQx4_ASAP7_75t_SL

MACRO DFFLQNx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFLQNx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 1.012 0.027 1.062 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx1_ASAP7_75t_SL

MACRO DFFLQNx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFLQNx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.115 0.243 ;
			RECT 1.097 0.027 1.115 0.243 ;
			RECT 1.012 0.027 1.115 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx2_ASAP7_75t_SL

MACRO DFFLQNx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFLQNx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.012 0.225 1.171 0.243 ;
			RECT 1.153 0.027 1.171 0.243 ;
			RECT 1.011 0.027 1.171 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.09 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQNx3_ASAP7_75t_SL

MACRO DFFLQx4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DFFLQx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.125 0.225 1.333 0.243 ;
			RECT 1.313 0.027 1.333 0.243 ;
			RECT 1.125 0.027 1.333 0.045 ;
			RECT 1.125 0.201 1.143 0.243 ;
			RECT 1.125 0.027 1.143 0.069 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.164 0.117 0.236 ;
			RECT 0.072 0.07 0.117 0.106 ;
			RECT 0.099 0.034 0.117 0.106 ;
			RECT 0.072 0.164 0.117 0.2 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.012 0.225 1.098 0.243 ;
			RECT 1.08 0.027 1.098 0.243 ;
			RECT 1.08 0.127 1.175 0.145 ;
			RECT 1.012 0.027 1.098 0.045 ;
			RECT 0.85 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.774 0.027 0.792 0.119 ;
			RECT 0.774 0.027 0.954 0.045 ;
			RECT 0.688 0.225 0.738 0.243 ;
			RECT 0.72 0.027 0.738 0.243 ;
			RECT 0.72 0.153 0.9 0.171 ;
			RECT 0.882 0.117 0.9 0.171 ;
			RECT 0.828 0.117 0.846 0.171 ;
			RECT 0.634 0.027 0.738 0.045 ;
			RECT 0.576 0.225 0.63 0.243 ;
			RECT 0.612 0.081 0.63 0.243 ;
			RECT 0.496 0.081 0.63 0.099 ;
			RECT 0.585 0.034 0.603 0.099 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.581 0.14 ;
			RECT 0.418 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.145 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.121 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.99 0.122 1.008 0.167 ;
			RECT 0.666 0.099 0.684 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.167 ;
			RECT 0.342 0.126 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.877 0.144 1.013 0.162 ;
			RECT 0.229 0.144 0.689 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			LAYER V1 ;
			RECT 0.99 0.144 1.008 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.15 0.18 0.168 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DFFLQx4_ASAP7_75t_SL

MACRO DHLx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DHLx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.742 0.027 0.792 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.72 0.122 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.743 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx1_ASAP7_75t_SL

MACRO DHLx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DHLx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.741 0.216 0.85 0.234 ;
			RECT 0.832 0.036 0.85 0.234 ;
			RECT 0.742 0.036 0.85 0.054 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.72 0.09 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.797 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx2_ASAP7_75t_SL

MACRO DHLx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DHLx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.918 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.688 0.225 0.9 0.243 ;
			RECT 0.882 0.027 0.9 0.243 ;
			RECT 0.688 0.027 0.9 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.918 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.918 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.096 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.121 0.581 0.139 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.106 0.36 0.207 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.18 0.198 0.198 ;
			RECT 0.18 0.126 0.198 0.198 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.828 0.09 0.846 0.167 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.72 0.09 0.738 0.167 ;
			RECT 0.504 0.164 0.522 0.207 ;
			RECT 0.396 0.106 0.414 0.171 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.851 0.162 ;
			RECT 0.019 0.18 0.527 0.198 ;
			RECT 0.229 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.153 0.18 0.171 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END DHLx3_ASAP7_75t_SL

MACRO DLLx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DLLx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.735 0.027 0.792 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.72 0.106 0.738 0.2 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.743 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.72 0.144 0.738 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx1_ASAP7_75t_SL

MACRO DLLx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DLLx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.688 0.225 0.847 0.243 ;
			RECT 0.829 0.027 0.847 0.243 ;
			RECT 0.688 0.027 0.847 0.045 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.8 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx2_ASAP7_75t_SL

MACRO DLLx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN DLLx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.918 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.742 0.216 0.901 0.234 ;
			RECT 0.882 0.036 0.901 0.234 ;
			RECT 0.742 0.036 0.901 0.054 ;

		END 

	END Q
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.153 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.117 ;
			RECT 0.099 0.034 0.117 0.117 ;
			RECT 0.072 0.153 0.117 0.189 ;
			RECT 0.072 0.081 0.09 0.189 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.325 0.243 ;
			RECT 0.288 0.027 0.325 0.045 ;
			RECT 0.288 0.027 0.306 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.918 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.918 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.58 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.504 0.027 0.522 0.097 ;
			RECT 0.504 0.027 0.63 0.045 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.45 0.122 0.58 0.14 ;
			RECT 0.414 0.027 0.468 0.045 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.148 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.138 0.126 0.198 0.144 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 0.774 0.09 0.792 0.167 ;
			RECT 0.504 0.165 0.522 0.203 ;
			RECT 0.396 0.106 0.414 0.2 ;
			RECT 0.342 0.106 0.36 0.203 ;
			LAYER M2 ;
			RECT 0.45 0.144 0.8 0.162 ;
			RECT 0.229 0.18 0.527 0.198 ;
			RECT 0.019 0.144 0.414 0.162 ;
			LAYER V1 ;
			RECT 0.774 0.144 0.792 0.162 ;
			RECT 0.504 0.18 0.522 0.198 ;
			RECT 0.45 0.144 0.468 0.162 ;
			RECT 0.396 0.144 0.414 0.162 ;
			RECT 0.342 0.18 0.36 0.198 ;
			RECT 0.234 0.18 0.252 0.198 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END DLLx3_ASAP7_75t_SL

MACRO FAx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN FAx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN CON
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.128 0.072 0.543 0.09 ;
			LAYER M1 ;
			RECT 0.515 0.072 0.543 0.09 ;
			RECT 0.504 0.09 0.533 0.108 ;
			RECT 0.504 0.09 0.522 0.149 ;
			RECT 0.124 0.072 0.282 0.09 ;
			RECT 0.124 0.189 0.23 0.207 ;
			RECT 0.124 0.072 0.142 0.207 ;
			LAYER V1 ;
			RECT 0.133 0.072 0.151 0.09 ;
			RECT 0.52 0.072 0.538 0.09 ;

		END 

	END CON
	PIN SN
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.324 0.225 0.495 0.243 ;
			RECT 0.477 0.184 0.495 0.243 ;
			RECT 0.477 0.027 0.495 0.068 ;
			RECT 0.324 0.027 0.495 0.045 ;
			RECT 0.324 0.027 0.342 0.243 ;

		END 

	END SN
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.059 0.18 0.627 0.198 ;
			LAYER M1 ;
			RECT 0.599 0.18 0.63 0.198 ;
			RECT 0.612 0.121 0.63 0.198 ;
			RECT 0.383 0.18 0.414 0.198 ;
			RECT 0.396 0.121 0.414 0.198 ;
			RECT 0.059 0.18 0.09 0.198 ;
			RECT 0.072 0.121 0.09 0.198 ;
			LAYER V1 ;
			RECT 0.064 0.18 0.082 0.198 ;
			RECT 0.388 0.18 0.406 0.198 ;
			RECT 0.604 0.18 0.622 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.167 0.144 0.689 0.162 ;
			LAYER M1 ;
			RECT 0.666 0.121 0.684 0.167 ;
			RECT 0.288 0.121 0.306 0.167 ;
			RECT 0.167 0.144 0.198 0.162 ;
			RECT 0.18 0.121 0.198 0.162 ;
			LAYER V1 ;
			RECT 0.172 0.144 0.19 0.162 ;
			RECT 0.288 0.144 0.306 0.162 ;
			RECT 0.666 0.144 0.684 0.162 ;

		END 

	END B
	PIN CI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.108 0.587 0.126 ;
			LAYER M1 ;
			RECT 0.558 0.108 0.587 0.126 ;
			RECT 0.558 0.108 0.576 0.149 ;
			RECT 0.45 0.103 0.468 0.149 ;
			RECT 0.226 0.108 0.263 0.126 ;
			RECT 0.234 0.108 0.252 0.149 ;
			LAYER V1 ;
			RECT 0.234 0.108 0.252 0.126 ;
			RECT 0.45 0.108 0.468 0.126 ;
			RECT 0.564 0.108 0.582 0.126 ;

		END 

	END CI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.027 0.662 0.045 ;
			RECT 0.526 0.225 0.662 0.243 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END FAx1_ASAP7_75t_SL

MACRO FILLER_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN FILLER_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.108 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.108 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.108 0.279 ;

		END 

	END VDD

END FILLER_ASAP7_75t_SL

MACRO FILLERxp5_ASAP7_75t_SL
	CLASS CORE SPACER ;
	FOREIGN FILLERxp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.054 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.054 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.054 0.279 ;

		END 

	END VDD

END FILLERxp5_ASAP7_75t_SL

MACRO HAxp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN HAxp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN CON
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.162 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.075 0.18 0.243 ;

		END 

	END CON
	PIN SN
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.423 0.027 0.468 0.045 ;

		END 

	END SN
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.15 ;
			RECT 0.207 0.063 0.36 0.081 ;
			RECT 0.207 0.027 0.225 0.081 ;
			RECT 0.018 0.027 0.225 0.045 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.027 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.106 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.387 0.045 ;

	END

END HAxp5_ASAP7_75t_SL

MACRO HB1xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN HB1xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.117 0.243 ;
			RECT 0.099 0.153 0.117 0.243 ;
			RECT 0.099 0.153 0.144 0.171 ;
			RECT 0.126 0.099 0.144 0.171 ;
			RECT 0.099 0.099 0.144 0.117 ;
			RECT 0.099 0.027 0.117 0.117 ;
			RECT 0.04 0.027 0.117 0.045 ;

	END

END HB1xp67_ASAP7_75t_SL

MACRO HB2xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN HB2xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.202 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.04 0.027 0.144 0.045 ;

	END

END HB2xp67_ASAP7_75t_SL

MACRO HB3xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN HB3xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.256 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.18 0.126 0.257 0.144 ;
			RECT 0.04 0.027 0.198 0.045 ;

	END

END HB3xp67_ASAP7_75t_SL

MACRO HB4xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN HB4xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.081 0.055 0.099 ;
			RECT 0.018 0.081 0.036 0.207 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.18 0.126 0.311 0.144 ;
			RECT 0.04 0.027 0.198 0.045 ;

	END

END HB4xp67_ASAP7_75t_SL

MACRO ICGx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.972 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.879 0.027 0.954 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.972 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.972 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx1_ASAP7_75t_SL

MACRO ICGx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.026 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 1.008 0.243 ;
			RECT 0.99 0.027 1.008 0.243 ;
			RECT 0.879 0.027 1.008 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.026 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.026 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx2_ASAP7_75t_SL

MACRO ICGx2p67DC_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx2p67DC_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx2p67DC_ASAP7_75t_SL

MACRO ICGx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.899 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.879 0.027 1.062 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx3_ASAP7_75t_SL

MACRO ICGx4DC_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx4DC_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx4DC_ASAP7_75t_SL

MACRO ICGx4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.134 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.89 0.225 1.062 0.243 ;
			RECT 1.044 0.027 1.062 0.243 ;
			RECT 0.889 0.027 1.062 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.134 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.134 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx4_ASAP7_75t_SL

MACRO ICGx5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.188 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.89 0.225 1.17 0.243 ;
			RECT 1.152 0.027 1.17 0.243 ;
			RECT 0.889 0.027 1.17 0.045 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.144 0.635 0.162 ;
			LAYER M1 ;
			RECT 0.612 0.178 0.765 0.196 ;
			RECT 0.747 0.142 0.765 0.196 ;
			RECT 0.612 0.116 0.63 0.196 ;
			RECT 0.396 0.144 0.447 0.162 ;
			RECT 0.396 0.12 0.414 0.162 ;
			RECT 0.234 0.119 0.252 0.184 ;
			LAYER V1 ;
			RECT 0.234 0.144 0.252 0.162 ;
			RECT 0.414 0.144 0.432 0.162 ;
			RECT 0.612 0.144 0.63 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.199 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.199 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.188 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.188 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.688 0.222 0.846 0.24 ;
			RECT 0.828 0.188 0.846 0.24 ;
			RECT 0.828 0.188 0.9 0.206 ;
			RECT 0.882 0.063 0.9 0.206 ;
			RECT 0.742 0.063 0.9 0.081 ;
			RECT 0.256 0.223 0.367 0.241 ;
			RECT 0.349 0.027 0.367 0.241 ;
			RECT 0.349 0.181 0.473 0.199 ;
			RECT 0.828 0.099 0.846 0.147 ;
			RECT 0.666 0.027 0.684 0.147 ;
			RECT 0.666 0.099 0.846 0.117 ;
			RECT 0.31 0.027 0.684 0.045 ;
			RECT 0.559 0.223 0.609 0.241 ;
			RECT 0.559 0.077 0.577 0.241 ;
			RECT 0.559 0.077 0.609 0.095 ;
			RECT 0.468 0.224 0.522 0.242 ;
			RECT 0.503 0.073 0.522 0.242 ;
			RECT 0.392 0.073 0.522 0.091 ;
			RECT 0.288 0.18 0.324 0.198 ;
			RECT 0.288 0.072 0.306 0.198 ;
			RECT 0.257 0.072 0.306 0.09 ;
			RECT 0.037 0.224 0.198 0.242 ;
			RECT 0.18 0.027 0.198 0.242 ;
			RECT 0.089 0.027 0.198 0.045 ;
			LAYER M2 ;
			RECT 0.296 0.18 0.582 0.198 ;
			LAYER V1 ;
			RECT 0.559 0.18 0.577 0.198 ;
			RECT 0.301 0.18 0.319 0.198 ;

	END

END ICGx5_ASAP7_75t_SL

MACRO ICGx5p33DC_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx5p33DC_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx5p33DC_ASAP7_75t_SL

MACRO ICGx6p67DC_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx6p67DC_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx6p67DC_ASAP7_75t_SL

MACRO ICGx8DC_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN ICGx8DC_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.592 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN GCLK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 2.465 0.225 2.52 0.243 ;
			RECT 2.502 0.027 2.52 0.243 ;
			RECT 2.445 0.027 2.52 0.045 ;
			RECT 1.925 0.225 1.98 0.243 ;
			RECT 1.962 0.027 1.98 0.243 ;
			RECT 1.905 0.027 1.98 0.045 ;
			RECT 0.612 0.027 0.687 0.045 ;
			RECT 0.612 0.225 0.667 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.072 0.027 0.147 0.045 ;
			RECT 0.072 0.225 0.127 0.243 ;
			RECT 0.072 0.027 0.09 0.243 ;
			LAYER M2 ;
			RECT 0.061 0.036 2.531 0.054 ;
			LAYER V1 ;
			RECT 0.072 0.036 0.09 0.054 ;
			RECT 0.612 0.036 0.63 0.054 ;
			RECT 1.962 0.036 1.98 0.054 ;
			RECT 2.502 0.036 2.52 0.054 ;

		END 

	END GCLK
	PIN CLK
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 2.281 0.171 2.35 0.189 ;
			RECT 2.332 0.135 2.35 0.189 ;
			RECT 2.292 0.135 2.35 0.153 ;
			RECT 1.638 0.178 1.791 0.196 ;
			RECT 1.773 0.142 1.791 0.196 ;
			RECT 1.638 0.116 1.656 0.196 ;
			RECT 1.422 0.144 1.473 0.162 ;
			RECT 1.422 0.12 1.44 0.162 ;
			RECT 1.26 0.119 1.278 0.184 ;
			RECT 0.801 0.178 0.954 0.196 ;
			RECT 0.936 0.116 0.954 0.196 ;
			RECT 0.801 0.142 0.819 0.196 ;
			RECT 0.248 0.171 0.317 0.189 ;
			RECT 0.248 0.135 0.306 0.153 ;
			RECT 0.248 0.135 0.266 0.189 ;
			LAYER M2 ;
			RECT 0.235 0.144 2.358 0.162 ;
			LAYER V1 ;
			RECT 0.248 0.144 0.266 0.162 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.44 0.144 1.458 0.162 ;
			RECT 1.638 0.144 1.656 0.162 ;
			RECT 2.332 0.144 2.35 0.162 ;

		END 

	END CLK
	PIN ENA
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.076 0.172 1.116 0.199 ;
			RECT 1.098 0.07 1.116 0.199 ;
			RECT 1.032 0.222 1.095 0.241 ;
			RECT 1.076 0.172 1.095 0.241 ;
			LAYER M2 ;
			RECT 0.982 0.216 1.237 0.234 ;
			LAYER V1 ;
			RECT 1.076 0.216 1.095 0.234 ;

		END 

	END ENA
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.152 0.07 1.17 0.199 ;
			LAYER M2 ;
			RECT 0.982 0.072 1.237 0.09 ;
			LAYER V1 ;
			RECT 1.152 0.072 1.17 0.09 ;

		END 

	END SE
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 2.592 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 2.592 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 2.254 0.222 2.412 0.24 ;
			RECT 2.394 0.188 2.412 0.24 ;
			RECT 2.394 0.188 2.466 0.206 ;
			RECT 2.448 0.063 2.466 0.206 ;
			RECT 2.308 0.063 2.466 0.081 ;
			RECT 2.394 0.099 2.412 0.147 ;
			RECT 2.232 0.099 2.25 0.147 ;
			RECT 2.232 0.099 2.412 0.117 ;
			RECT 2.124 0.126 2.18 0.144 ;
			RECT 2.124 0.09 2.142 0.144 ;
			RECT 2.038 0.09 2.19 0.108 ;
			RECT 2.019 0.162 2.174 0.18 ;
			RECT 2.07 0.126 2.088 0.18 ;
			RECT 2.03 0.126 2.088 0.144 ;
			RECT 1.714 0.222 1.872 0.24 ;
			RECT 1.854 0.188 1.872 0.24 ;
			RECT 1.854 0.188 1.926 0.206 ;
			RECT 1.908 0.063 1.926 0.206 ;
			RECT 1.768 0.063 1.926 0.081 ;
			RECT 1.282 0.223 1.393 0.241 ;
			RECT 1.375 0.027 1.393 0.241 ;
			RECT 1.375 0.181 1.499 0.199 ;
			RECT 1.854 0.099 1.872 0.147 ;
			RECT 1.692 0.027 1.71 0.147 ;
			RECT 1.692 0.099 1.872 0.117 ;
			RECT 1.336 0.027 1.71 0.045 ;
			RECT 1.585 0.223 1.635 0.241 ;
			RECT 1.585 0.077 1.603 0.241 ;
			RECT 1.585 0.077 1.635 0.095 ;
			RECT 1.494 0.224 1.548 0.242 ;
			RECT 1.529 0.073 1.548 0.242 ;
			RECT 1.418 0.073 1.548 0.091 ;
			RECT 1.314 0.18 1.35 0.198 ;
			RECT 1.314 0.072 1.332 0.198 ;
			RECT 1.283 0.072 1.332 0.09 ;
			RECT 1.12 0.224 1.224 0.242 ;
			RECT 1.206 0.027 1.224 0.242 ;
			RECT 1.115 0.027 1.224 0.045 ;
			RECT 0.957 0.223 1.007 0.241 ;
			RECT 0.989 0.077 1.007 0.241 ;
			RECT 0.957 0.077 1.007 0.095 ;
			RECT 0.882 0.099 0.9 0.147 ;
			RECT 0.72 0.099 0.738 0.147 ;
			RECT 0.72 0.099 0.9 0.117 ;
			RECT 0.72 0.222 0.878 0.24 ;
			RECT 0.72 0.188 0.738 0.24 ;
			RECT 0.666 0.188 0.738 0.206 ;
			RECT 0.666 0.063 0.684 0.206 ;
			RECT 0.666 0.063 0.824 0.081 ;
			RECT 0.418 0.162 0.573 0.18 ;
			RECT 0.504 0.126 0.522 0.18 ;
			RECT 0.504 0.126 0.562 0.144 ;
			RECT 0.412 0.126 0.468 0.144 ;
			RECT 0.45 0.09 0.468 0.144 ;
			RECT 0.402 0.09 0.554 0.108 ;
			RECT 0.342 0.099 0.36 0.147 ;
			RECT 0.18 0.099 0.198 0.147 ;
			RECT 0.18 0.099 0.36 0.117 ;
			RECT 0.18 0.222 0.338 0.24 ;
			RECT 0.18 0.188 0.198 0.24 ;
			RECT 0.126 0.188 0.198 0.206 ;
			RECT 0.126 0.063 0.144 0.206 ;
			RECT 0.126 0.063 0.284 0.081 ;
			LAYER M2 ;
			RECT 0.336 0.108 2.256 0.126 ;
			RECT 0.982 0.18 1.608 0.198 ;
			LAYER V1 ;
			RECT 2.232 0.108 2.25 0.126 ;
			RECT 1.692 0.108 1.71 0.126 ;
			RECT 1.585 0.18 1.603 0.198 ;
			RECT 1.327 0.18 1.345 0.198 ;
			RECT 0.989 0.18 1.007 0.198 ;
			RECT 0.882 0.108 0.9 0.126 ;
			RECT 0.342 0.108 0.36 0.126 ;

	END

END ICGx8DC_ASAP7_75t_SL

MACRO INVx11_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx11_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.684 0.243 ;
			RECT 0.666 0.027 0.684 0.243 ;
			RECT 0.094 0.027 0.684 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD

END INVx11_ASAP7_75t_SL

MACRO INVx13_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx13_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.094 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD

END INVx13_ASAP7_75t_SL

MACRO INVx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVx1_ASAP7_75t_SL

MACRO INVx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END INVx2_ASAP7_75t_SL

MACRO INVx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.252 0.243 ;
			RECT 0.234 0.027 0.252 0.243 ;
			RECT 0.094 0.027 0.252 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END INVx3_ASAP7_75t_SL

MACRO INVx4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END INVx4_ASAP7_75t_SL

MACRO INVx5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.094 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END INVx5_ASAP7_75t_SL

MACRO INVx6_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx6_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.094 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD

END INVx6_ASAP7_75t_SL

MACRO INVx8_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVx8_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.522 0.243 ;
			RECT 0.504 0.027 0.522 0.243 ;
			RECT 0.094 0.027 0.522 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD

END INVx8_ASAP7_75t_SL

MACRO INVxp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVxp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVxp33_ASAP7_75t_SL

MACRO INVxp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN INVxp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.027 0.144 0.243 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END INVxp67_ASAP7_75t_SL

MACRO MAJIxp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN MAJIxp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.255 0.189 0.361 0.207 ;
			RECT 0.343 0.063 0.361 0.207 ;
			RECT 0.255 0.063 0.361 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.126 0.257 0.144 ;
			RECT 0.018 0.189 0.198 0.207 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.027 0.338 0.045 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END MAJIxp5_ASAP7_75t_SL

MACRO MAJx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN MAJx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.364 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.333 0.207 ;
			RECT 0.315 0.106 0.333 0.207 ;
			RECT 0.283 0.126 0.333 0.144 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.121 0.126 0.198 0.144 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.063 0.036 0.207 ;
			RECT 0.368 0.063 0.386 0.149 ;
			RECT 0.018 0.063 0.386 0.081 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END MAJx2_ASAP7_75t_SL

MACRO MAJx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN MAJx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.504 0.243 ;
			RECT 0.364 0.027 0.504 0.045 ;
			RECT 0.45 0.027 0.468 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.189 0.333 0.207 ;
			RECT 0.315 0.106 0.333 0.207 ;
			RECT 0.283 0.126 0.333 0.144 ;
			RECT 0.18 0.126 0.198 0.207 ;
			RECT 0.121 0.126 0.198 0.144 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.189 0.123 0.207 ;
			RECT 0.018 0.063 0.036 0.207 ;
			RECT 0.368 0.063 0.386 0.149 ;
			RECT 0.018 0.063 0.386 0.081 ;
			RECT 0.04 0.027 0.284 0.045 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END MAJx3_ASAP7_75t_SL

MACRO NAND2x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND2x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.202 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.065 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END NAND2x1_ASAP7_75t_SL

MACRO NAND2x1p5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND2x1p5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.261 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.063 0.338 0.081 ;
			RECT 0.094 0.027 0.225 0.045 ;

	END

END NAND2x1p5_ASAP7_75t_SL

MACRO NAND2x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND2x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.418 0.063 0.522 0.081 ;
			RECT 0.018 0.063 0.122 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.242 0.189 0.279 0.207 ;
			RECT 0.261 0.106 0.279 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.177 ;
			RECT 0.322 0.099 0.468 0.117 ;
			RECT 0.322 0.063 0.34 0.117 ;
			RECT 0.2 0.063 0.34 0.081 ;
			RECT 0.072 0.099 0.218 0.117 ;
			RECT 0.2 0.063 0.218 0.117 ;
			RECT 0.072 0.189 0.109 0.207 ;
			RECT 0.072 0.099 0.09 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.5 0.045 ;

	END

END NAND2x2_ASAP7_75t_SL

MACRO NAND2xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND2xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.143 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NAND2xp33_ASAP7_75t_SL

MACRO NAND2xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND2xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.143 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.106 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NAND2xp5_ASAP7_75t_SL

MACRO NAND2xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND2xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.202 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.125 0.095 0.143 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.063 0.055 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.106 0.252 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END NAND2xp67_ASAP7_75t_SL

MACRO NAND3x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND3x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.418 0.063 0.576 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.402 0.18 0.468 0.198 ;
			RECT 0.45 0.108 0.468 0.198 ;
			RECT 0.4 0.108 0.468 0.126 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.243 0.18 0.306 0.198 ;
			RECT 0.288 0.108 0.306 0.198 ;
			RECT 0.246 0.108 0.306 0.126 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.061 0.103 0.079 0.203 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.5 0.045 ;
			RECT 0.094 0.063 0.338 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END NAND3x1_ASAP7_75t_SL

MACRO NAND3x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND3x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 1.062 0.243 ;
			RECT 1.044 0.063 1.062 0.243 ;
			RECT 0.904 0.063 1.062 0.081 ;
			RECT 0.018 0.063 0.176 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.169 0.18 0.908 0.198 ;
			LAYER M1 ;
			RECT 0.866 0.189 0.903 0.207 ;
			RECT 0.885 0.108 0.903 0.207 ;
			RECT 0.174 0.189 0.211 0.207 ;
			RECT 0.174 0.106 0.192 0.207 ;
			LAYER V1 ;
			RECT 0.174 0.18 0.192 0.198 ;
			RECT 0.885 0.18 0.903 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.338 0.189 0.743 0.207 ;
			RECT 0.725 0.106 0.743 0.207 ;
			RECT 0.338 0.106 0.356 0.207 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.547 0.106 0.565 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.742 0.027 0.986 0.045 ;
			RECT 0.256 0.063 0.824 0.081 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.094 0.027 0.338 0.045 ;

	END

END NAND3x2_ASAP7_75t_SL

MACRO NAND3xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND3xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END NAND3xp33_ASAP7_75t_SL

MACRO NAND4xp25_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND4xp25_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.256 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.034 0.09 0.2 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END NAND4xp25_ASAP7_75t_SL

MACRO NAND4xp75_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND4xp75_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.738 0.243 ;
			RECT 0.72 0.063 0.738 0.243 ;
			RECT 0.58 0.063 0.738 0.081 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.106 0.63 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.101 0.549 0.119 ;
			RECT 0.531 0.07 0.549 0.119 ;
			RECT 0.504 0.101 0.522 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.101 0.306 0.2 ;
			RECT 0.207 0.101 0.306 0.119 ;
			RECT 0.207 0.07 0.225 0.119 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.057 0.243 ;
			RECT 0.018 0.027 0.057 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.412 0.027 0.666 0.045 ;
			RECT 0.256 0.063 0.499 0.081 ;
			RECT 0.092 0.027 0.34 0.045 ;

	END

END NAND4xp75_ASAP7_75t_SL

MACRO NAND5xp2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NAND5xp2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.009 0.225 0.317 0.243 ;
			RECT 0.009 0.027 0.07 0.045 ;
			RECT 0.009 0.027 0.027 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.034 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.034 0.198 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.034 0.252 0.2 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.034 0.306 0.2 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END NAND5xp2_ASAP7_75t_SL

MACRO NOR2x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR2x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.23 0.144 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END NOR2x1_ASAP7_75t_SL

MACRO NOR2x1p5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR2x1p5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.094 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.084 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.063 0.163 0.081 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.189 0.338 0.207 ;
			RECT 0.094 0.225 0.225 0.243 ;

	END

END NOR2x1p5_ASAP7_75t_SL

MACRO NOR2x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR2x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.189 0.522 0.207 ;
			RECT 0.504 0.027 0.522 0.207 ;
			RECT 0.018 0.027 0.522 0.045 ;
			RECT 0.018 0.189 0.122 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.063 0.279 0.164 ;
			RECT 0.242 0.063 0.279 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.322 0.153 0.468 0.171 ;
			RECT 0.45 0.093 0.468 0.171 ;
			RECT 0.2 0.189 0.34 0.207 ;
			RECT 0.322 0.153 0.34 0.207 ;
			RECT 0.2 0.153 0.218 0.207 ;
			RECT 0.072 0.153 0.218 0.171 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.5 0.243 ;

	END

END NOR2x2_ASAP7_75t_SL

MACRO NOR2xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR2xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.216 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.143 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.094 0.027 0.198 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.225 0.055 0.243 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.216 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.216 0.279 ;

		END 

	END VDD

END NOR2xp33_ASAP7_75t_SL

MACRO NOR2xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR2xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.189 0.306 0.207 ;
			RECT 0.288 0.027 0.306 0.207 ;
			RECT 0.148 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.127 0.095 0.145 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.257 0.144 ;
			RECT 0.126 0.063 0.163 0.081 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END NOR2xp67_ASAP7_75t_SL

MACRO NOR3x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR3x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.418 0.189 0.576 0.207 ;
			RECT 0.558 0.027 0.576 0.207 ;
			RECT 0.202 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.153 0.468 0.171 ;
			RECT 0.45 0.063 0.468 0.171 ;
			RECT 0.396 0.063 0.468 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.153 0.306 0.171 ;
			RECT 0.288 0.063 0.306 0.171 ;
			RECT 0.234 0.063 0.306 0.081 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.189 0.055 0.207 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.225 0.5 0.243 ;
			RECT 0.094 0.189 0.338 0.207 ;
			RECT 0.04 0.225 0.176 0.243 ;

	END

END NOR3x1_ASAP7_75t_SL

MACRO NOR3x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR3x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.08 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.904 0.189 1.062 0.207 ;
			RECT 1.044 0.027 1.062 0.207 ;
			RECT 0.018 0.027 1.062 0.045 ;
			RECT 0.018 0.189 0.176 0.207 ;
			RECT 0.018 0.027 0.036 0.207 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.169 0.072 0.908 0.09 ;
			LAYER M1 ;
			RECT 0.885 0.063 0.903 0.162 ;
			RECT 0.866 0.063 0.903 0.081 ;
			RECT 0.174 0.063 0.211 0.081 ;
			RECT 0.174 0.063 0.192 0.164 ;
			LAYER V1 ;
			RECT 0.174 0.072 0.192 0.09 ;
			RECT 0.885 0.072 0.903 0.09 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.725 0.063 0.743 0.164 ;
			RECT 0.338 0.063 0.743 0.081 ;
			RECT 0.338 0.063 0.356 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.547 0.106 0.565 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.08 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.08 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.742 0.225 0.986 0.243 ;
			RECT 0.256 0.189 0.824 0.207 ;
			RECT 0.418 0.225 0.662 0.243 ;
			RECT 0.094 0.225 0.338 0.243 ;

	END

END NOR3x2_ASAP7_75t_SL

MACRO NOR3xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR3xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.176 0.045 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD

END NOR3xp33_ASAP7_75t_SL

MACRO NOR4xp25_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR4xp25_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.04 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD

END NOR4xp25_ASAP7_75t_SL

MACRO NOR4xp75_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR4xp75_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.756 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.58 0.189 0.738 0.207 ;
			RECT 0.72 0.027 0.738 0.207 ;
			RECT 0.094 0.027 0.738 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.07 0.63 0.164 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.531 0.151 0.549 0.2 ;
			RECT 0.504 0.151 0.549 0.169 ;
			RECT 0.504 0.07 0.522 0.169 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.151 0.306 0.169 ;
			RECT 0.288 0.07 0.306 0.169 ;
			RECT 0.207 0.151 0.225 0.2 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.225 0.057 0.243 ;
			RECT 0.018 0.027 0.057 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.756 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.756 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.412 0.225 0.666 0.243 ;
			RECT 0.256 0.189 0.499 0.207 ;
			RECT 0.092 0.225 0.34 0.243 ;

	END

END NOR4xp75_ASAP7_75t_SL

MACRO NOR5xp2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN NOR5xp2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.017 0.027 0.338 0.045 ;
			RECT 0.017 0.225 0.07 0.243 ;
			RECT 0.017 0.027 0.037 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD

END NOR5xp2_ASAP7_75t_SL

MACRO O2A1O1Ixp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN O2A1O1Ixp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.094 0.027 0.306 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.206 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.225 0.243 ;
			RECT 0.04 0.063 0.176 0.081 ;

	END

END O2A1O1Ixp33_ASAP7_75t_SL

MACRO O2A1O1Ixp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN O2A1O1Ixp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.315 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.063 0.252 0.164 ;
			RECT 0.072 0.063 0.252 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.164 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.164 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.189 0.338 0.207 ;
			RECT 0.148 0.027 0.279 0.045 ;
			RECT 0.094 0.225 0.23 0.243 ;

	END

END O2A1O1Ixp5_ASAP7_75t_SL

MACRO OA211x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA211x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.296 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.286 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.164 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.252 0.243 ;
			RECT 0.234 0.189 0.252 0.243 ;
			RECT 0.234 0.189 0.306 0.207 ;
			RECT 0.288 0.063 0.306 0.207 ;
			RECT 0.099 0.063 0.306 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OA211x2_ASAP7_75t_SL

MACRO OA21x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA21x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.256 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.153 0.239 0.171 ;
			RECT 0.18 0.106 0.198 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.225 0.224 0.243 ;
			RECT 0.206 0.189 0.224 0.243 ;
			RECT 0.206 0.189 0.306 0.207 ;
			RECT 0.288 0.063 0.306 0.207 ;
			RECT 0.099 0.063 0.306 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OA21x2_ASAP7_75t_SL

MACRO OA221x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA221x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.864 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.225 0.117 0.243 ;
			RECT 0.099 0.189 0.117 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.215 0.189 0.252 0.207 ;
			RECT 0.234 0.099 0.252 0.207 ;
			RECT 0.215 0.099 0.252 0.117 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.189 0.379 0.207 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.593 0.189 0.63 0.207 ;
			RECT 0.612 0.099 0.63 0.207 ;
			RECT 0.593 0.099 0.63 0.117 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.099 0.522 0.207 ;
			RECT 0.485 0.099 0.522 0.117 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.72 0.189 0.757 0.207 ;
			RECT 0.72 0.099 0.757 0.117 ;
			RECT 0.72 0.099 0.738 0.207 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.864 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.864 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.144 0.225 0.846 0.243 ;
			RECT 0.828 0.063 0.846 0.243 ;
			RECT 0.144 0.126 0.162 0.243 ;
			RECT 0.121 0.126 0.162 0.144 ;
			RECT 0.741 0.063 0.846 0.081 ;
			RECT 0.472 0.027 0.824 0.045 ;
			RECT 0.202 0.063 0.668 0.081 ;

	END

END OA221x2_ASAP7_75t_SL

MACRO OA222x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA222x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.531 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.526 0.027 0.63 0.045 ;
			RECT 0.531 0.189 0.549 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.009 0.225 0.504 0.243 ;
			RECT 0.486 0.126 0.504 0.243 ;
			RECT 0.009 0.063 0.027 0.243 ;
			RECT 0.486 0.126 0.554 0.144 ;
			RECT 0.009 0.063 0.122 0.081 ;
			RECT 0.202 0.063 0.36 0.081 ;
			RECT 0.342 0.027 0.36 0.081 ;
			RECT 0.342 0.027 0.468 0.045 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OA222x2_ASAP7_75t_SL

MACRO OA22x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA22x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.071 0.225 0.122 0.243 ;
			RECT 0.071 0.027 0.122 0.045 ;
			RECT 0.071 0.027 0.091 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.236 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.063 0.414 0.2 ;
			RECT 0.367 0.063 0.414 0.081 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.18 0.225 0.392 0.243 ;
			RECT 0.18 0.063 0.198 0.243 ;
			RECT 0.137 0.126 0.198 0.144 ;
			RECT 0.18 0.063 0.333 0.081 ;
			RECT 0.256 0.027 0.5 0.045 ;

	END

END OA22x2_ASAP7_75t_SL

MACRO OA31x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA31x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.81 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.225 0.792 0.243 ;
			RECT 0.774 0.027 0.792 0.243 ;
			RECT 0.693 0.027 0.792 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.053 0.189 0.09 0.207 ;
			RECT 0.072 0.099 0.09 0.207 ;
			RECT 0.053 0.099 0.09 0.117 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.126 0.189 0.163 0.207 ;
			RECT 0.126 0.106 0.144 0.207 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.126 0.414 0.144 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.323 0.063 0.36 0.081 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.153 0.522 0.171 ;
			RECT 0.504 0.106 0.522 0.171 ;

		END 

	END B1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.81 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.81 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.369 0.189 0.576 0.207 ;
			RECT 0.558 0.063 0.576 0.207 ;
			RECT 0.558 0.126 0.667 0.144 ;
			RECT 0.418 0.063 0.576 0.081 ;
			RECT 0.317 0.225 0.446 0.243 ;
			RECT 0.317 0.189 0.335 0.243 ;
			RECT 0.202 0.189 0.335 0.207 ;
			RECT 0.094 0.027 0.5 0.045 ;
			RECT 0.04 0.063 0.284 0.081 ;
			RECT 0.04 0.225 0.284 0.243 ;

	END

END OA31x2_ASAP7_75t_SL

MACRO OA331x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA331x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.166 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.099 0.186 0.117 0.243 ;
			RECT 0.072 0.186 0.117 0.204 ;
			RECT 0.072 0.115 0.09 0.204 ;
			RECT 0.471 0.063 0.522 0.081 ;
			RECT 0.234 0.063 0.393 0.081 ;
			RECT 0.234 0.027 0.252 0.081 ;
			RECT 0.148 0.027 0.252 0.045 ;
			RECT 0.308 0.027 0.447 0.045 ;

	END

END OA331x1_ASAP7_75t_SL

MACRO OA331x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA331x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.045 0.225 0.122 0.243 ;
			RECT 0.045 0.027 0.122 0.045 ;
			RECT 0.045 0.027 0.063 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.166 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.153 0.186 0.171 0.243 ;
			RECT 0.126 0.186 0.171 0.204 ;
			RECT 0.126 0.115 0.144 0.204 ;
			RECT 0.525 0.063 0.576 0.081 ;
			RECT 0.288 0.063 0.447 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.202 0.027 0.306 0.045 ;
			RECT 0.362 0.027 0.501 0.045 ;

	END

END OA331x2_ASAP7_75t_SL

MACRO OA332x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA332x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.094 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.126 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.126 0.189 0.144 0.243 ;
			RECT 0.072 0.189 0.144 0.207 ;
			RECT 0.072 0.119 0.09 0.207 ;
			RECT 0.471 0.063 0.576 0.081 ;
			RECT 0.234 0.063 0.393 0.081 ;
			RECT 0.234 0.027 0.252 0.081 ;
			RECT 0.146 0.027 0.252 0.045 ;
			RECT 0.308 0.027 0.556 0.045 ;

	END

END OA332x1_ASAP7_75t_SL

MACRO OA332x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA332x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.137 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.18 0.225 0.63 0.243 ;
			RECT 0.612 0.063 0.63 0.243 ;
			RECT 0.18 0.189 0.198 0.243 ;
			RECT 0.126 0.189 0.198 0.207 ;
			RECT 0.126 0.119 0.144 0.207 ;
			RECT 0.525 0.063 0.63 0.081 ;
			RECT 0.288 0.063 0.447 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.2 0.027 0.306 0.045 ;
			RECT 0.362 0.027 0.61 0.045 ;

	END

END OA332x2_ASAP7_75t_SL

MACRO OA333x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA333x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.225 0.63 0.243 ;
			RECT 0.612 0.063 0.63 0.243 ;
			RECT 0.099 0.186 0.117 0.243 ;
			RECT 0.072 0.186 0.117 0.204 ;
			RECT 0.072 0.115 0.09 0.204 ;
			RECT 0.467 0.063 0.63 0.081 ;
			RECT 0.232 0.063 0.394 0.081 ;
			RECT 0.232 0.027 0.25 0.081 ;
			RECT 0.147 0.027 0.25 0.045 ;
			RECT 0.309 0.027 0.569 0.045 ;

	END

END OA333x1_ASAP7_75t_SL

MACRO OA333x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA333x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.225 0.122 0.243 ;
			RECT 0.072 0.027 0.122 0.045 ;
			RECT 0.072 0.027 0.09 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.612 0.106 0.63 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.558 0.106 0.576 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.164 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.153 0.225 0.684 0.243 ;
			RECT 0.666 0.063 0.684 0.243 ;
			RECT 0.153 0.186 0.171 0.243 ;
			RECT 0.126 0.186 0.171 0.204 ;
			RECT 0.126 0.115 0.144 0.204 ;
			RECT 0.521 0.063 0.684 0.081 ;
			RECT 0.286 0.063 0.448 0.081 ;
			RECT 0.286 0.027 0.304 0.081 ;
			RECT 0.201 0.027 0.304 0.045 ;
			RECT 0.363 0.027 0.623 0.045 ;

	END

END OA333x2_ASAP7_75t_SL

MACRO OA33x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OA33x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.225 0.117 0.243 ;
			RECT 0.099 0.189 0.117 0.243 ;
			RECT 0.062 0.189 0.117 0.207 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.144 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.144 0.126 0.162 0.243 ;
			RECT 0.121 0.126 0.162 0.144 ;
			RECT 0.364 0.063 0.522 0.081 ;
			RECT 0.202 0.027 0.446 0.045 ;

	END

END OA33x2_ASAP7_75t_SL

MACRO OAI211xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI211xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.099 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.09 0.144 ;
			RECT 0.018 0.07 0.036 0.2 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI211xp5_ASAP7_75t_SL

MACRO OAI21x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI21x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.369 0.027 0.414 0.045 ;
			RECT 0.018 0.027 0.063 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.189 0.306 0.207 ;
			RECT 0.288 0.106 0.306 0.207 ;
			RECT 0.126 0.106 0.144 0.207 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.19 0.127 0.256 0.145 ;
			RECT 0.19 0.099 0.227 0.171 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.072 0.063 0.36 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.027 0.333 0.045 ;

	END

END OAI21x1_ASAP7_75t_SL

MACRO OAI21xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI21xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.099 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.203 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI21xp33_ASAP7_75t_SL

MACRO OAI21xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI21xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.27 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.148 0.225 0.252 0.243 ;
			RECT 0.234 0.063 0.252 0.243 ;
			RECT 0.099 0.063 0.252 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.203 ;

		END 

	END A2
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.171 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.27 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.27 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI21xp5_ASAP7_75t_SL

MACRO OAI221xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI221xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.23 0.243 ;
			RECT 0.018 0.063 0.123 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.201 0.063 0.339 0.081 ;
			RECT 0.04 0.027 0.176 0.045 ;

	END

END OAI221xp5_ASAP7_75t_SL

MACRO OAI222xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI222xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.522 0.243 ;
			RECT 0.504 0.055 0.522 0.243 ;
			RECT 0.018 0.063 0.122 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.07 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.07 0.468 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.063 0.36 0.081 ;
			RECT 0.342 0.027 0.36 0.081 ;
			RECT 0.342 0.027 0.468 0.045 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI222xp33_ASAP7_75t_SL

MACRO OAI22x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI22x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.038 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.309 0.063 0.522 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.153 0.379 0.171 ;
			RECT 0.342 0.099 0.379 0.117 ;
			RECT 0.342 0.099 0.36 0.171 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.189 0.468 0.207 ;
			RECT 0.45 0.099 0.468 0.207 ;
			RECT 0.431 0.099 0.468 0.117 ;
			RECT 0.288 0.118 0.306 0.207 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.161 0.153 0.198 0.171 ;
			RECT 0.18 0.063 0.198 0.171 ;
			RECT 0.161 0.063 0.198 0.081 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.189 0.252 0.207 ;
			RECT 0.234 0.116 0.252 0.207 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.207 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.5 0.045 ;

	END

END OAI22x1_ASAP7_75t_SL

MACRO OAI22xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI22xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.063 0.117 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.225 0.275 0.243 ;
			RECT 0.234 0.07 0.252 0.243 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI22xp33_ASAP7_75t_SL

MACRO OAI22xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI22xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.176 0.243 ;
			RECT 0.018 0.063 0.117 0.081 ;
			RECT 0.018 0.063 0.036 0.243 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END A2
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.225 0.275 0.243 ;
			RECT 0.234 0.07 0.252 0.243 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.063 0.198 0.164 ;
			RECT 0.151 0.063 0.198 0.081 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.027 0.284 0.045 ;

	END

END OAI22xp5_ASAP7_75t_SL

MACRO OAI311xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI311xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.198 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.31 0.027 0.36 0.045 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.2 ;

		END 

	END B1
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.027 0.234 0.045 ;

	END

END OAI311xp33_ASAP7_75t_SL

MACRO OAI31xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI31xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.306 0.243 ;
			RECT 0.288 0.063 0.306 0.243 ;
			RECT 0.256 0.063 0.306 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.093 0.027 0.23 0.045 ;

	END

END OAI31xp33_ASAP7_75t_SL

MACRO OAI31xp67_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI31xp67_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.702 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.202 0.063 0.663 0.081 ;
			RECT 0.202 0.189 0.252 0.207 ;
			RECT 0.234 0.063 0.252 0.207 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.666 0.126 0.684 0.198 ;
			RECT 0.553 0.126 0.684 0.144 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.126 0.419 0.144 ;
			RECT 0.288 0.126 0.306 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.07 0.036 0.236 ;

		END 

	END A3
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.126 0.203 0.144 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.702 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.702 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.526 0.225 0.663 0.243 ;
			RECT 0.364 0.189 0.608 0.207 ;
			RECT 0.04 0.027 0.554 0.045 ;
			RECT 0.094 0.225 0.446 0.243 ;

	END

END OAI31xp67_ASAP7_75t_SL

MACRO OAI321xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI321xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.198 0.225 0.414 0.243 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.31 0.063 0.414 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.095 0.144 ;
			RECT 0.018 0.034 0.036 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B2
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.256 0.027 0.396 0.045 ;
			RECT 0.094 0.063 0.23 0.081 ;

	END

END OAI321xp33_ASAP7_75t_SL

MACRO OAI322xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI322xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.147 0.225 0.468 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.364 0.063 0.468 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.105 0.306 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END B2
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.105 0.36 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.202 0.027 0.45 0.045 ;
			RECT 0.039 0.063 0.284 0.081 ;

	END

END OAI322xp33_ASAP7_75t_SL

MACRO OAI32xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI32xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.04 0.225 0.36 0.243 ;
			RECT 0.342 0.063 0.36 0.243 ;
			RECT 0.256 0.063 0.36 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.063 0.222 0.081 ;
			RECT 0.18 0.063 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.099 0.027 0.338 0.045 ;

	END

END OAI32xp33_ASAP7_75t_SL

MACRO OAI331xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI331xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.468 0.243 ;
			RECT 0.45 0.063 0.468 0.243 ;
			RECT 0.417 0.063 0.468 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C1
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.393 0.045 ;
			RECT 0.092 0.063 0.339 0.081 ;

	END

END OAI331xp33_ASAP7_75t_SL

MACRO OAI332xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI332xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.54 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.522 0.243 ;
			RECT 0.504 0.063 0.522 0.243 ;
			RECT 0.417 0.063 0.522 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END C2
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.54 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.54 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.502 0.045 ;
			RECT 0.092 0.063 0.339 0.081 ;

	END

END OAI332xp33_ASAP7_75t_SL

MACRO OAI333xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI333xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.576 0.243 ;
			RECT 0.558 0.063 0.576 0.243 ;
			RECT 0.413 0.063 0.576 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.504 0.106 0.522 0.2 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.106 0.468 0.2 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.2 ;

		END 

	END C1
	PIN C2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END C2
	PIN C3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END C3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.254 0.027 0.515 0.045 ;
			RECT 0.094 0.063 0.34 0.081 ;

	END

END OAI333xp33_ASAP7_75t_SL

MACRO OAI33xp33_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OAI33xp33_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.201 0.225 0.414 0.243 ;
			RECT 0.396 0.063 0.414 0.243 ;
			RECT 0.256 0.063 0.414 0.081 ;

		END 

	END Y
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.236 ;

		END 

	END A1
	PIN A2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END A2
	PIN A3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END A3
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.106 0.252 0.2 ;

		END 

	END B1
	PIN B2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.2 ;

		END 

	END B2
	PIN B3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.106 0.36 0.2 ;

		END 

	END B3
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.092 0.027 0.338 0.045 ;

	END

END OAI33xp33_ASAP7_75t_SL

MACRO OR2x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR2x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.306 0.243 ;
			RECT 0.288 0.027 0.306 0.243 ;
			RECT 0.207 0.027 0.306 0.045 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.077 0.144 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.186 0.243 ;
			RECT 0.168 0.027 0.186 0.243 ;
			RECT 0.168 0.126 0.227 0.144 ;
			RECT 0.094 0.027 0.186 0.045 ;

	END

END OR2x2_ASAP7_75t_SL

MACRO OR2x4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR2x4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.207 0.027 0.414 0.045 ;
			RECT 0.315 0.184 0.333 0.243 ;
			RECT 0.315 0.027 0.333 0.086 ;
			RECT 0.207 0.184 0.225 0.243 ;
			RECT 0.207 0.027 0.225 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.126 0.077 0.144 ;
			RECT 0.018 0.027 0.055 0.045 ;
			RECT 0.018 0.027 0.036 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.187 0.243 ;
			RECT 0.169 0.027 0.187 0.243 ;
			RECT 0.169 0.126 0.227 0.144 ;
			RECT 0.094 0.027 0.187 0.045 ;

	END

END OR2x4_ASAP7_75t_SL

MACRO OR2x6_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR2x6_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.225 0.63 0.243 ;
			RECT 0.612 0.027 0.63 0.243 ;
			RECT 0.31 0.027 0.63 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.063 0.144 0.122 ;
			RECT 0.018 0.063 0.144 0.081 ;
			RECT 0.018 0.063 0.036 0.236 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.153 0.252 0.171 ;
			RECT 0.234 0.121 0.252 0.171 ;
			RECT 0.072 0.106 0.09 0.236 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.148 0.189 0.306 0.207 ;
			RECT 0.288 0.07 0.306 0.207 ;
			RECT 0.234 0.07 0.306 0.088 ;
			RECT 0.234 0.027 0.252 0.088 ;
			RECT 0.094 0.027 0.252 0.045 ;

	END

END OR2x6_ASAP7_75t_SL

MACRO OR3x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR3x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.324 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.183 0.306 0.201 ;
			RECT 0.288 0.076 0.306 0.201 ;
			RECT 0.261 0.076 0.306 0.094 ;
			RECT 0.261 0.183 0.279 0.235 ;
			RECT 0.261 0.034 0.279 0.094 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.324 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.324 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.234 0.243 ;
			RECT 0.216 0.027 0.234 0.243 ;
			RECT 0.216 0.126 0.262 0.144 ;
			RECT 0.04 0.027 0.234 0.045 ;

	END

END OR3x1_ASAP7_75t_SL

MACRO OR3x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR3x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.261 0.027 0.36 0.045 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.24 0.243 ;
			RECT 0.222 0.027 0.24 0.243 ;
			RECT 0.222 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.24 0.045 ;

	END

END OR3x2_ASAP7_75t_SL

MACRO OR3x4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR3x4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.261 0.027 0.468 0.045 ;
			RECT 0.369 0.184 0.387 0.243 ;
			RECT 0.369 0.027 0.387 0.086 ;
			RECT 0.261 0.184 0.279 0.243 ;
			RECT 0.261 0.027 0.279 0.086 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.2 ;

		END 

	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.04 0.225 0.241 0.243 ;
			RECT 0.223 0.027 0.241 0.243 ;
			RECT 0.223 0.126 0.284 0.144 ;
			RECT 0.04 0.027 0.241 0.045 ;

	END

END OR3x4_ASAP7_75t_SL

MACRO OR4x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR4x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.378 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.027 0.068 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.106 0.144 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.378 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.378 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.072 0.066 0.09 0.152 ;
			RECT 0.072 0.066 0.117 0.084 ;
			RECT 0.099 0.027 0.117 0.084 ;
			RECT 0.099 0.027 0.36 0.045 ;

	END

END OR4x1_ASAP7_75t_SL

MACRO OR4x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR4x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.018 0.225 0.122 0.243 ;
			RECT 0.018 0.027 0.122 0.045 ;
			RECT 0.018 0.027 0.036 0.243 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.07 0.36 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.07 0.306 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.106 0.198 0.236 ;

		END 

	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.364 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.099 0.063 0.117 0.149 ;
			RECT 0.099 0.063 0.171 0.081 ;
			RECT 0.153 0.027 0.171 0.081 ;
			RECT 0.153 0.027 0.414 0.045 ;

	END

END OR4x2_ASAP7_75t_SL

MACRO OR5x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR5x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.432 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.35 0.225 0.414 0.243 ;
			RECT 0.396 0.027 0.414 0.243 ;
			RECT 0.349 0.027 0.414 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.432 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.432 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.07 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.288 0.063 0.36 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.018 0.027 0.306 0.045 ;

	END

END OR5x1_ASAP7_75t_SL

MACRO OR5x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN OR5x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.364 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.343 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.07 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.236 ;

		END 

	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.18 0.07 0.198 0.236 ;

		END 

	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.234 0.07 0.252 0.236 ;

		END 

	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.288 0.106 0.306 0.236 ;

		END 

	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.07 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.342 0.063 0.36 0.154 ;
			RECT 0.288 0.063 0.36 0.081 ;
			RECT 0.288 0.027 0.306 0.081 ;
			RECT 0.018 0.027 0.306 0.045 ;

	END

END OR5x2_ASAP7_75t_SL

MACRO SDFHx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFHx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.332 0.243 ;
			RECT 1.314 0.027 1.332 0.243 ;
			RECT 1.282 0.027 1.332 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.099 0.185 0.117 0.236 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.185 0.117 0.203 ;
			RECT 0.072 0.081 0.09 0.203 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.284 0.108 0.436 0.126 ;
			LAYER M1 ;
			RECT 0.396 0.106 0.414 0.164 ;
			LAYER V1 ;
			RECT 0.396 0.108 0.414 0.126 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.467 0.108 0.59 0.126 ;
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;
			LAYER V1 ;
			RECT 0.504 0.108 0.522 0.126 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.797 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.021 0.225 0.068 0.243 ;
			RECT 0.021 0.027 0.039 0.243 ;
			RECT 0.021 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.016 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.021 0.144 0.039 0.162 ;

	END

END SDFHx1_ASAP7_75t_SL

MACRO SDFHx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFHx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.282 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.019 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx2_ASAP7_75t_SL

MACRO SDFHx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFHx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.458 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.44 0.243 ;
			RECT 1.422 0.027 1.44 0.243 ;
			RECT 1.282 0.027 1.44 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.458 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.458 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			RECT 0.126 0.121 0.144 0.167 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.019 0.144 0.9 0.162 ;
			RECT 0.175 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.18 0.198 0.198 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx3_ASAP7_75t_SL

MACRO SDFHx4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFHx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.674 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.444 0.225 1.656 0.243 ;
			RECT 1.637 0.027 1.656 0.243 ;
			RECT 1.444 0.027 1.656 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.164 ;
			RECT 0.378 0.225 0.459 0.243 ;
			RECT 0.378 0.099 0.468 0.117 ;
			RECT 0.378 0.099 0.396 0.243 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.599 0.081 ;
			RECT 0.558 0.063 0.576 0.164 ;
			RECT 0.234 0.126 0.289 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;
			LAYER V1 ;
			RECT 0.234 0.072 0.252 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.027 0.767 0.045 ;
			RECT 0.639 0.063 0.711 0.081 ;
			RECT 0.693 0.027 0.711 0.081 ;
			RECT 0.612 0.106 0.657 0.124 ;
			RECT 0.639 0.063 0.657 0.124 ;
			RECT 0.612 0.106 0.63 0.164 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.674 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.674 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.059 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.368 0.126 1.447 0.144 ;
			RECT 1.242 0.126 1.283 0.144 ;
			RECT 1.242 0.027 1.26 0.144 ;
			RECT 1.113 0.027 1.386 0.045 ;
			RECT 1.206 0.182 1.332 0.2 ;
			RECT 1.314 0.081 1.332 0.2 ;
			RECT 1.206 0.106 1.224 0.2 ;
			RECT 1.287 0.081 1.332 0.099 ;
			RECT 0.882 0.063 0.9 0.164 ;
			RECT 0.882 0.063 0.981 0.081 ;
			RECT 0.801 0.225 0.954 0.243 ;
			RECT 0.936 0.106 0.954 0.243 ;
			RECT 0.801 0.189 0.819 0.243 ;
			RECT 0.738 0.189 0.819 0.207 ;
			RECT 0.738 0.07 0.756 0.207 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.504 0.063 0.522 0.164 ;
			RECT 0.342 0.063 0.522 0.081 ;
			RECT 0.31 0.027 0.36 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.126 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.144 0.047 0.162 ;
			RECT 0.009 0.027 0.09 0.045 ;
			RECT 1.152 0.106 1.17 0.2 ;
			RECT 1.098 0.07 1.116 0.164 ;
			RECT 1.044 0.106 1.062 0.2 ;
			RECT 0.828 0.07 0.846 0.167 ;
			RECT 0.774 0.07 0.792 0.164 ;
			RECT 0.58 0.225 0.77 0.243 ;
			RECT 0.684 0.121 0.702 0.167 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.423 0.189 0.662 0.207 ;
			RECT 0.126 0.106 0.144 0.2 ;
			LAYER M2 ;
			RECT 0.019 0.144 1.175 0.162 ;
			RECT 0.175 0.108 1.121 0.126 ;
			LAYER V1 ;
			RECT 1.152 0.144 1.17 0.162 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 1.044 0.144 1.062 0.162 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.108 0.792 0.126 ;
			RECT 0.684 0.144 0.702 0.162 ;
			RECT 0.18 0.108 0.198 0.126 ;
			RECT 0.126 0.144 0.144 0.162 ;
			RECT 0.024 0.144 0.042 0.162 ;

	END

END SDFHx4_ASAP7_75t_SL

MACRO SDFLx1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFLx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.35 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.332 0.243 ;
			RECT 1.314 0.027 1.332 0.243 ;
			RECT 1.282 0.027 1.332 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.35 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.35 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.797 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx1_ASAP7_75t_SL

MACRO SDFLx2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFLx2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.404 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.282 0.027 1.386 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.404 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.404 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx2_ASAP7_75t_SL

MACRO SDFLx3_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFLx3_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.458 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.282 0.225 1.44 0.243 ;
			RECT 1.422 0.027 1.44 0.243 ;
			RECT 1.282 0.027 1.44 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.081 0.117 0.099 ;
			RECT 0.099 0.034 0.117 0.099 ;
			RECT 0.072 0.081 0.09 0.164 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.396 0.099 0.433 0.117 ;
			RECT 0.396 0.099 0.414 0.164 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.211 0.036 1.229 0.054 ;
			LAYER M1 ;
			RECT 1.206 0.027 1.25 0.045 ;
			RECT 1.206 0.027 1.224 0.2 ;
			RECT 0.216 0.126 0.311 0.144 ;
			RECT 0.216 0.027 0.258 0.045 ;
			RECT 0.216 0.027 0.234 0.144 ;
			LAYER V1 ;
			RECT 0.216 0.036 0.234 0.054 ;
			RECT 1.206 0.036 1.224 0.054 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.485 0.189 0.522 0.207 ;
			RECT 0.504 0.106 0.522 0.207 ;
			RECT 0.461 0.126 0.522 0.144 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.458 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.458 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.152 0.225 1.202 0.243 ;
			RECT 1.152 0.034 1.17 0.243 ;
			RECT 1.066 0.225 1.116 0.243 ;
			RECT 1.098 0.027 1.116 0.243 ;
			RECT 0.99 0.027 1.008 0.119 ;
			RECT 0.99 0.027 1.116 0.045 ;
			RECT 0.904 0.225 0.954 0.243 ;
			RECT 0.936 0.027 0.954 0.243 ;
			RECT 0.936 0.153 1.062 0.171 ;
			RECT 1.044 0.117 1.062 0.171 ;
			RECT 0.85 0.027 0.954 0.045 ;
			RECT 0.792 0.225 0.846 0.243 ;
			RECT 0.828 0.081 0.846 0.243 ;
			RECT 0.72 0.081 0.846 0.099 ;
			RECT 0.801 0.045 0.819 0.099 ;
			RECT 0.72 0.062 0.738 0.099 ;
			RECT 0.58 0.225 0.702 0.243 ;
			RECT 0.684 0.027 0.702 0.243 ;
			RECT 0.684 0.122 0.792 0.14 ;
			RECT 0.634 0.027 0.702 0.045 ;
			RECT 0.612 0.153 0.649 0.171 ;
			RECT 0.612 0.106 0.63 0.171 ;
			RECT 0.558 0.189 0.595 0.207 ;
			RECT 0.558 0.106 0.576 0.207 ;
			RECT 0.261 0.081 0.306 0.099 ;
			RECT 0.288 0.027 0.306 0.099 ;
			RECT 0.288 0.027 0.5 0.045 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.342 0.063 0.379 0.081 ;
			RECT 0.126 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.148 0.027 0.198 0.045 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.18 0.047 0.198 ;
			RECT 0.009 0.027 0.068 0.045 ;
			RECT 1.26 0.09 1.278 0.2 ;
			RECT 0.882 0.101 0.9 0.167 ;
			RECT 0.72 0.165 0.738 0.207 ;
			RECT 0.418 0.063 0.609 0.081 ;
			RECT 0.255 0.225 0.5 0.243 ;
			RECT 0.309 0.189 0.447 0.207 ;
			LAYER M2 ;
			RECT 0.936 0.144 1.283 0.162 ;
			RECT 0.337 0.072 1.175 0.09 ;
			RECT 0.175 0.144 0.9 0.162 ;
			RECT 0.019 0.18 0.743 0.198 ;
			LAYER V1 ;
			RECT 1.26 0.144 1.278 0.162 ;
			RECT 1.152 0.072 1.17 0.09 ;
			RECT 0.936 0.144 0.954 0.162 ;
			RECT 0.882 0.144 0.9 0.162 ;
			RECT 0.72 0.18 0.738 0.198 ;
			RECT 0.612 0.144 0.63 0.162 ;
			RECT 0.558 0.18 0.576 0.198 ;
			RECT 0.342 0.072 0.36 0.09 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.024 0.18 0.042 0.198 ;

	END

END SDFLx3_ASAP7_75t_SL

MACRO SDFLx4_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN SDFLx4_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.674 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER M1 ;
			RECT 1.444 0.225 1.656 0.243 ;
			RECT 1.637 0.027 1.656 0.243 ;
			RECT 1.444 0.027 1.656 0.045 ;

		END 

	END QN
	PIN CLK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER M1 ;
			RECT 0.072 0.063 0.109 0.081 ;
			RECT 0.072 0.063 0.09 0.2 ;

		END 

	END CLK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.45 0.099 0.468 0.164 ;
			RECT 0.378 0.225 0.459 0.243 ;
			RECT 0.378 0.099 0.468 0.117 ;
			RECT 0.378 0.099 0.396 0.243 ;

		END 

	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER M2 ;
			RECT 0.229 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.599 0.081 ;
			RECT 0.558 0.063 0.576 0.164 ;
			RECT 0.234 0.126 0.289 0.144 ;
			RECT 0.234 0.225 0.271 0.243 ;
			RECT 0.234 0.027 0.271 0.045 ;
			RECT 0.234 0.027 0.252 0.243 ;
			LAYER V1 ;
			RECT 0.234 0.072 0.252 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER M1 ;
			RECT 0.693 0.027 0.767 0.045 ;
			RECT 0.639 0.063 0.711 0.081 ;
			RECT 0.693 0.027 0.711 0.081 ;
			RECT 0.612 0.106 0.657 0.124 ;
			RECT 0.639 0.063 0.657 0.124 ;
			RECT 0.612 0.106 0.63 0.164 ;

		END 

	END SI
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 1.674 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 1.674 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 1.059 0.225 1.386 0.243 ;
			RECT 1.368 0.027 1.386 0.243 ;
			RECT 1.368 0.126 1.447 0.144 ;
			RECT 1.242 0.126 1.283 0.144 ;
			RECT 1.242 0.027 1.26 0.144 ;
			RECT 1.113 0.027 1.386 0.045 ;
			RECT 1.206 0.182 1.332 0.2 ;
			RECT 1.314 0.081 1.332 0.2 ;
			RECT 1.206 0.106 1.224 0.2 ;
			RECT 1.287 0.081 1.332 0.099 ;
			RECT 0.882 0.063 0.9 0.164 ;
			RECT 0.882 0.063 0.981 0.081 ;
			RECT 0.801 0.225 0.954 0.243 ;
			RECT 0.936 0.106 0.954 0.243 ;
			RECT 0.801 0.189 0.819 0.243 ;
			RECT 0.738 0.189 0.819 0.207 ;
			RECT 0.738 0.07 0.756 0.207 ;
			RECT 0.31 0.225 0.36 0.243 ;
			RECT 0.342 0.027 0.36 0.243 ;
			RECT 0.504 0.063 0.522 0.164 ;
			RECT 0.342 0.063 0.522 0.081 ;
			RECT 0.31 0.027 0.36 0.045 ;
			RECT 0.148 0.225 0.198 0.243 ;
			RECT 0.18 0.027 0.198 0.243 ;
			RECT 0.126 0.027 0.198 0.045 ;
			RECT 0.009 0.225 0.068 0.243 ;
			RECT 0.009 0.027 0.027 0.243 ;
			RECT 0.009 0.108 0.047 0.126 ;
			RECT 0.009 0.027 0.09 0.045 ;
			RECT 1.152 0.106 1.17 0.2 ;
			RECT 1.098 0.07 1.116 0.164 ;
			RECT 1.044 0.106 1.062 0.2 ;
			RECT 0.828 0.07 0.846 0.167 ;
			RECT 0.774 0.07 0.792 0.164 ;
			RECT 0.58 0.225 0.77 0.243 ;
			RECT 0.684 0.121 0.702 0.167 ;
			RECT 0.418 0.027 0.662 0.045 ;
			RECT 0.423 0.189 0.662 0.207 ;
			RECT 0.126 0.103 0.144 0.2 ;
			LAYER M2 ;
			RECT 0.175 0.144 1.175 0.162 ;
			RECT 0.019 0.108 1.121 0.126 ;
			LAYER V1 ;
			RECT 1.152 0.144 1.17 0.162 ;
			RECT 1.098 0.108 1.116 0.126 ;
			RECT 1.044 0.144 1.062 0.162 ;
			RECT 0.828 0.144 0.846 0.162 ;
			RECT 0.774 0.108 0.792 0.126 ;
			RECT 0.684 0.144 0.702 0.162 ;
			RECT 0.18 0.144 0.198 0.162 ;
			RECT 0.126 0.108 0.144 0.126 ;
			RECT 0.024 0.108 0.042 0.126 ;

	END

END SDFLx4_ASAP7_75t_SL

MACRO TAPCELL_ASAP7_75t_SL
	CLASS CORE WELLTAP ;
	FOREIGN TAPCELL_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.108 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.108 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.108 0.279 ;

		END 

	END VDD

END TAPCELL_ASAP7_75t_SL

MACRO TAPCELL_WITH_FILLER_ASAP7_75t_SL
	CLASS CORE WELLTAP ;
	FOREIGN TAPCELL_WITH_FILLER_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD

END TAPCELL_WITH_FILLER_ASAP7_75t_SL

MACRO TIEHIx1_ASAP7_75t_SL
	CLASS CORE TIEHIGH ;
	FOREIGN TIEHIx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN H
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.094 0.225 0.144 0.243 ;
			RECT 0.126 0.07 0.144 0.243 ;
			RECT 0.067 0.07 0.144 0.088 ;

		END 

	END H
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.155 0.095 0.173 ;
			RECT 0.018 0.027 0.036 0.173 ;
			RECT 0.018 0.027 0.068 0.045 ;

	END

END TIEHIx1_ASAP7_75t_SL

MACRO TIELOx1_ASAP7_75t_SL
	CLASS CORE TIELOW ;
	FOREIGN TIELOx1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.162 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN L
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.067 0.182 0.144 0.2 ;
			RECT 0.126 0.027 0.144 0.2 ;
			RECT 0.094 0.027 0.144 0.045 ;

		END 

	END L
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.162 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.162 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.068 0.243 ;
			RECT 0.018 0.097 0.036 0.243 ;
			RECT 0.018 0.097 0.095 0.115 ;

	END

END TIELOx1_ASAP7_75t_SL

MACRO XNOR2x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN XNOR2x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.612 0.243 ;
			RECT 0.45 0.077 0.468 0.243 ;
			RECT 0.418 0.077 0.468 0.095 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.121 0.18 0.581 0.198 ;
			LAYER M1 ;
			RECT 0.526 0.189 0.576 0.207 ;
			RECT 0.558 0.121 0.576 0.207 ;
			RECT 0.107 0.189 0.144 0.207 ;
			RECT 0.126 0.121 0.144 0.207 ;
			LAYER V1 ;
			RECT 0.126 0.18 0.144 0.198 ;
			RECT 0.558 0.18 0.576 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.298 0.072 0.527 0.09 ;
			LAYER M1 ;
			RECT 0.504 0.07 0.522 0.152 ;
			RECT 0.305 0.126 0.365 0.144 ;
			RECT 0.305 0.067 0.323 0.144 ;
			RECT 0.213 0.067 0.323 0.085 ;
			RECT 0.213 0.027 0.231 0.085 ;
			RECT 0.018 0.027 0.231 0.045 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.027 0.036 0.236 ;
			LAYER V1 ;
			RECT 0.305 0.072 0.323 0.09 ;
			RECT 0.504 0.072 0.522 0.09 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.092 0.225 0.193 0.243 ;
			RECT 0.174 0.189 0.193 0.243 ;
			RECT 0.174 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.174 0.082 0.192 0.243 ;
			RECT 0.256 0.027 0.608 0.045 ;

	END

END XNOR2x1_ASAP7_75t_SL

MACRO XNOR2x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN XNOR2x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.472 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.261 0.225 0.44 0.243 ;
			RECT 0.422 0.126 0.44 0.243 ;
			RECT 0.391 0.126 0.44 0.144 ;
			RECT 0.261 0.183 0.279 0.243 ;
			RECT 0.126 0.183 0.279 0.201 ;
			RECT 0.126 0.12 0.144 0.201 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.189 0.38 0.207 ;
			RECT 0.342 0.107 0.36 0.207 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.063 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.477 0.063 0.495 0.151 ;
			RECT 0.423 0.063 0.495 0.081 ;
			RECT 0.423 0.027 0.441 0.081 ;
			RECT 0.018 0.027 0.441 0.045 ;
			RECT 0.302 0.063 0.32 0.195 ;
			RECT 0.072 0.063 0.09 0.149 ;
			RECT 0.072 0.063 0.392 0.081 ;
			RECT 0.099 0.225 0.23 0.243 ;

	END

END XNOR2x2_ASAP7_75t_SL

MACRO XNOR2xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN XNOR2xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.423 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.36 0.164 ;
			RECT 0.207 0.063 0.36 0.081 ;
			RECT 0.207 0.027 0.225 0.081 ;
			RECT 0.072 0.027 0.225 0.045 ;
			RECT 0.072 0.027 0.09 0.2 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.126 0.07 0.144 0.2 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.094 0.225 0.18 0.243 ;
			RECT 0.162 0.075 0.18 0.243 ;
			RECT 0.162 0.189 0.414 0.207 ;
			RECT 0.396 0.121 0.414 0.207 ;
			RECT 0.261 0.027 0.387 0.045 ;

	END

END XNOR2xp5_ASAP7_75t_SL

MACRO XOR2x1_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN XOR2x1_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.648 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.256 0.027 0.612 0.045 ;
			RECT 0.418 0.175 0.468 0.193 ;
			RECT 0.45 0.027 0.468 0.193 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.298 0.18 0.527 0.198 ;
			LAYER M1 ;
			RECT 0.504 0.118 0.522 0.2 ;
			RECT 0.305 0.126 0.365 0.144 ;
			RECT 0.213 0.185 0.323 0.203 ;
			RECT 0.305 0.126 0.323 0.203 ;
			RECT 0.018 0.225 0.231 0.243 ;
			RECT 0.213 0.185 0.231 0.243 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.243 ;
			LAYER V1 ;
			RECT 0.305 0.18 0.323 0.198 ;
			RECT 0.504 0.18 0.522 0.198 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M2 ;
			RECT 0.121 0.072 0.581 0.09 ;
			LAYER M1 ;
			RECT 0.558 0.063 0.576 0.149 ;
			RECT 0.526 0.063 0.576 0.081 ;
			RECT 0.126 0.063 0.144 0.149 ;
			RECT 0.107 0.063 0.144 0.081 ;
			LAYER V1 ;
			RECT 0.126 0.072 0.144 0.09 ;
			RECT 0.558 0.072 0.576 0.09 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.648 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.648 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.174 0.027 0.192 0.188 ;
			RECT 0.396 0.063 0.414 0.149 ;
			RECT 0.174 0.063 0.414 0.081 ;
			RECT 0.174 0.027 0.193 0.081 ;
			RECT 0.092 0.027 0.193 0.045 ;
			RECT 0.256 0.225 0.608 0.243 ;

	END

END XOR2x1_ASAP7_75t_SL

MACRO XOR2x2_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN XOR2x2_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.594 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.472 0.225 0.576 0.243 ;
			RECT 0.558 0.027 0.576 0.243 ;
			RECT 0.472 0.027 0.576 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.342 0.063 0.38 0.081 ;
			RECT 0.342 0.063 0.36 0.163 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.422 0.027 0.44 0.163 ;
			RECT 0.391 0.126 0.44 0.144 ;
			RECT 0.261 0.027 0.44 0.045 ;
			RECT 0.126 0.069 0.279 0.087 ;
			RECT 0.261 0.027 0.279 0.087 ;
			RECT 0.126 0.069 0.144 0.15 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.594 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.594 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.018 0.225 0.441 0.243 ;
			RECT 0.423 0.189 0.441 0.243 ;
			RECT 0.018 0.027 0.036 0.243 ;
			RECT 0.423 0.189 0.495 0.207 ;
			RECT 0.477 0.119 0.495 0.207 ;
			RECT 0.018 0.027 0.063 0.045 ;
			RECT 0.072 0.189 0.392 0.207 ;
			RECT 0.302 0.075 0.32 0.207 ;
			RECT 0.072 0.121 0.09 0.207 ;
			RECT 0.099 0.027 0.23 0.045 ;

	END

END XOR2x2_ASAP7_75t_SL

MACRO XOR2xp5_ASAP7_75t_SL
	CLASS CORE ;
	FOREIGN XOR2xp5_ASAP7_75t_SL 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.486 BY 0.27 ;
	SYMMETRY X Y ;
	SITE asap7sc7p5t ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.423 0.225 0.468 0.243 ;
			RECT 0.45 0.027 0.468 0.243 ;
			RECT 0.256 0.027 0.468 0.045 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.207 0.189 0.36 0.207 ;
			RECT 0.342 0.12 0.36 0.207 ;
			RECT 0.018 0.225 0.225 0.243 ;
			RECT 0.207 0.189 0.225 0.243 ;
			RECT 0.018 0.126 0.078 0.144 ;
			RECT 0.018 0.034 0.036 0.243 ;

		END 

	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 0.106 0.189 0.144 0.207 ;
			RECT 0.126 0.063 0.144 0.207 ;
			RECT 0.107 0.063 0.144 0.081 ;

		END 

	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 -0.009 0.486 0.009 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M1 ;
			RECT 0.0 0.261 0.486 0.279 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.162 0.027 0.18 0.195 ;
			RECT 0.396 0.063 0.414 0.149 ;
			RECT 0.162 0.063 0.414 0.081 ;
			RECT 0.094 0.027 0.18 0.045 ;
			RECT 0.256 0.225 0.387 0.243 ;

	END

END XOR2xp5_ASAP7_75t_SL

MACRO sram_asap7_16x256_1rw
	CLASS BLOCK ;
	FOREIGN sram_asap7_16x256_1rw 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 8.36 BY 16.8 ;
	SYMMETRY X Y ;
	PIN clk
		DIRECTION INPUT ;
		USE CLOCK ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.168 0.024 15.192 ;

		END 

	END clk
	PIN rd_out[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.808 0.024 5.832 ;

		END 

	END rd_out[15]
	PIN rd_out[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.424 0.024 5.448 ;

		END 

	END rd_out[14]
	PIN rd_out[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.04 0.024 5.064 ;

		END 

	END rd_out[13]
	PIN rd_out[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.656 0.024 4.68 ;

		END 

	END rd_out[12]
	PIN rd_out[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.272 0.024 4.296 ;

		END 

	END rd_out[11]
	PIN rd_out[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.888 0.024 3.912 ;

		END 

	END rd_out[10]
	PIN rd_out[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.504 0.024 3.528 ;

		END 

	END rd_out[9]
	PIN rd_out[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.12 0.024 3.144 ;

		END 

	END rd_out[8]
	PIN rd_out[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.736 0.024 2.76 ;

		END 

	END rd_out[7]
	PIN rd_out[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.352 0.024 2.376 ;

		END 

	END rd_out[6]
	PIN rd_out[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.968 0.024 1.992 ;

		END 

	END rd_out[5]
	PIN rd_out[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.584 0.024 1.608 ;

		END 

	END rd_out[4]
	PIN rd_out[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.2 0.024 1.224 ;

		END 

	END rd_out[3]
	PIN rd_out[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.816 0.024 0.84 ;

		END 

	END rd_out[2]
	PIN rd_out[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.432 0.024 0.456 ;

		END 

	END rd_out[1]
	PIN rd_out[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.048 0.024 0.072 ;

		END 

	END rd_out[0]
	PIN we_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.4 0.024 14.424 ;

		END 

	END we_in
	PIN ce_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.784 0.024 14.808 ;

		END 

	END ce_in
	PIN addr_in[7]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.352 0.024 14.376 ;

		END 

	END addr_in[7]
	PIN addr_in[6]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.968 0.024 13.992 ;

		END 

	END addr_in[6]
	PIN addr_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.584 0.024 13.608 ;

		END 

	END addr_in[5]
	PIN addr_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.2 0.024 13.224 ;

		END 

	END addr_in[4]
	PIN addr_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.816 0.024 12.84 ;

		END 

	END addr_in[3]
	PIN addr_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.432 0.024 12.456 ;

		END 

	END addr_in[2]
	PIN addr_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.048 0.024 12.072 ;

		END 

	END addr_in[1]
	PIN addr_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.664 0.024 11.688 ;

		END 

	END addr_in[0]
	PIN wd_in[15]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.616 0.024 11.64 ;

		END 

	END wd_in[15]
	PIN wd_in[14]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.232 0.024 11.256 ;

		END 

	END wd_in[14]
	PIN wd_in[13]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.848 0.024 10.872 ;

		END 

	END wd_in[13]
	PIN wd_in[12]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.464 0.024 10.488 ;

		END 

	END wd_in[12]
	PIN wd_in[11]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.08 0.024 10.104 ;

		END 

	END wd_in[11]
	PIN wd_in[10]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.696 0.024 9.72 ;

		END 

	END wd_in[10]
	PIN wd_in[9]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.312 0.024 9.336 ;

		END 

	END wd_in[9]
	PIN wd_in[8]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.928 0.024 8.952 ;

		END 

	END wd_in[8]
	PIN wd_in[7]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.544 0.024 8.568 ;

		END 

	END wd_in[7]
	PIN wd_in[6]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.16 0.024 8.184 ;

		END 

	END wd_in[6]
	PIN wd_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.776 0.024 7.8 ;

		END 

	END wd_in[5]
	PIN wd_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.392 0.024 7.416 ;

		END 

	END wd_in[4]
	PIN wd_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.008 0.024 7.032 ;

		END 

	END wd_in[3]
	PIN wd_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.624 0.024 6.648 ;

		END 

	END wd_in[2]
	PIN wd_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.24 0.024 6.264 ;

		END 

	END wd_in[1]
	PIN wd_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.856 0.024 5.88 ;

		END 

	END wd_in[0]
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.0 8.312 0.096 ;
			RECT 0.048 0.768 8.312 0.864 ;
			RECT 0.048 1.536 8.312 1.632 ;
			RECT 0.048 2.304 8.312 2.4 ;
			RECT 0.048 3.072 8.312 3.168 ;
			RECT 0.048 3.84 8.312 3.936 ;
			RECT 0.048 4.608 8.312 4.704 ;
			RECT 0.048 5.376 8.312 5.472 ;
			RECT 0.048 6.144 8.312 6.24 ;
			RECT 0.048 6.912 8.312 7.008 ;
			RECT 0.048 7.68 8.312 7.776 ;
			RECT 0.048 8.448 8.312 8.544 ;
			RECT 0.048 9.216 8.312 9.312 ;
			RECT 0.048 9.984 8.312 10.08 ;
			RECT 0.048 10.752 8.312 10.848 ;
			RECT 0.048 11.52 8.312 11.616 ;
			RECT 0.048 12.288 8.312 12.384 ;
			RECT 0.048 13.056 8.312 13.152 ;
			RECT 0.048 13.824 8.312 13.92 ;
			RECT 0.048 14.592 8.312 14.688 ;
			RECT 0.048 15.36 8.312 15.456 ;
			RECT 0.048 16.128 8.312 16.224 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.384 8.312 0.48 ;
			RECT 0.048 1.152 8.312 1.248 ;
			RECT 0.048 1.92 8.312 2.016 ;
			RECT 0.048 2.688 8.312 2.784 ;
			RECT 0.048 3.456 8.312 3.552 ;
			RECT 0.048 4.224 8.312 4.32 ;
			RECT 0.048 4.992 8.312 5.088 ;
			RECT 0.048 5.76 8.312 5.856 ;
			RECT 0.048 6.528 8.312 6.624 ;
			RECT 0.048 7.296 8.312 7.392 ;
			RECT 0.048 8.064 8.312 8.16 ;
			RECT 0.048 8.832 8.312 8.928 ;
			RECT 0.048 9.6 8.312 9.696 ;
			RECT 0.048 10.368 8.312 10.464 ;
			RECT 0.048 11.136 8.312 11.232 ;
			RECT 0.048 11.904 8.312 12.0 ;
			RECT 0.048 12.672 8.312 12.768 ;
			RECT 0.048 13.44 8.312 13.536 ;
			RECT 0.048 14.208 8.312 14.304 ;
			RECT 0.048 14.976 8.312 15.072 ;
			RECT 0.048 15.744 8.312 15.84 ;
			RECT 0.048 16.512 8.312 16.608 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.0 0.0 8.36 16.8 ;
			LAYER M2 ;
			RECT 0.0 0.0 8.36 16.8 ;
			LAYER M3 ;
			RECT 0.0 0.0 8.36 16.8 ;
			LAYER M4 ;
			RECT 0.024 0.0 0.048 16.8 ;
			RECT 8.312 0.0 8.36 16.8 ;
			RECT 0.048 0.0 8.312 0.0 ;
			RECT 0.048 0.096 8.312 0.384 ;
			RECT 0.048 0.48 8.312 0.768 ;
			RECT 0.048 0.864 8.312 1.152 ;
			RECT 0.048 1.248 8.312 1.536 ;
			RECT 0.048 1.632 8.312 1.92 ;
			RECT 0.048 2.016 8.312 2.304 ;
			RECT 0.048 2.4 8.312 2.688 ;
			RECT 0.048 2.784 8.312 3.072 ;
			RECT 0.048 3.168 8.312 3.456 ;
			RECT 0.048 3.552 8.312 3.84 ;
			RECT 0.048 3.936 8.312 4.224 ;
			RECT 0.048 4.32 8.312 4.608 ;
			RECT 0.048 4.704 8.312 4.992 ;
			RECT 0.048 5.088 8.312 5.376 ;
			RECT 0.048 5.472 8.312 5.76 ;
			RECT 0.048 5.856 8.312 6.144 ;
			RECT 0.048 6.24 8.312 6.528 ;
			RECT 0.048 6.624 8.312 6.912 ;
			RECT 0.048 7.008 8.312 7.296 ;
			RECT 0.048 7.392 8.312 7.68 ;
			RECT 0.048 7.776 8.312 8.064 ;
			RECT 0.048 8.16 8.312 8.448 ;
			RECT 0.048 8.544 8.312 8.832 ;
			RECT 0.048 8.928 8.312 9.216 ;
			RECT 0.048 9.312 8.312 9.6 ;
			RECT 0.048 9.696 8.312 9.984 ;
			RECT 0.048 10.08 8.312 10.368 ;
			RECT 0.048 10.464 8.312 10.752 ;
			RECT 0.048 10.848 8.312 11.136 ;
			RECT 0.048 11.232 8.312 11.52 ;
			RECT 0.048 11.616 8.312 11.904 ;
			RECT 0.048 12.0 8.312 12.288 ;
			RECT 0.048 12.384 8.312 12.672 ;
			RECT 0.048 12.768 8.312 13.056 ;
			RECT 0.048 13.152 8.312 13.44 ;
			RECT 0.048 13.536 8.312 13.824 ;
			RECT 0.048 13.92 8.312 14.208 ;
			RECT 0.048 14.304 8.312 14.592 ;
			RECT 0.048 14.688 8.312 14.976 ;
			RECT 0.048 15.072 8.312 15.36 ;
			RECT 0.048 15.456 8.312 15.744 ;
			RECT 0.048 15.84 8.312 16.128 ;
			RECT 0.048 16.224 8.312 16.512 ;
			RECT 0.048 16.608 8.312 16.8 ;
			RECT 0.0 0.0 0.024 0.048 ;
			RECT 0.0 0.072 0.024 0.432 ;
			RECT 0.0 0.456 0.024 0.816 ;
			RECT 0.0 0.84 0.024 1.2 ;
			RECT 0.0 1.224 0.024 1.584 ;
			RECT 0.0 1.608 0.024 1.968 ;
			RECT 0.0 1.992 0.024 2.352 ;
			RECT 0.0 2.376 0.024 2.736 ;
			RECT 0.0 2.76 0.024 3.12 ;
			RECT 0.0 3.144 0.024 3.504 ;
			RECT 0.0 3.528 0.024 3.888 ;
			RECT 0.0 3.912 0.024 4.272 ;
			RECT 0.0 4.296 0.024 4.656 ;
			RECT 0.0 4.68 0.024 5.04 ;
			RECT 0.0 5.064 0.024 5.424 ;
			RECT 0.0 5.448 0.024 5.808 ;
			RECT 0.0 5.832 0.024 5.856 ;
			RECT 0.0 5.88 0.024 6.24 ;
			RECT 0.0 6.264 0.024 6.624 ;
			RECT 0.0 6.648 0.024 7.008 ;
			RECT 0.0 7.032 0.024 7.392 ;
			RECT 0.0 7.416 0.024 7.776 ;
			RECT 0.0 7.8 0.024 8.16 ;
			RECT 0.0 8.184 0.024 8.544 ;
			RECT 0.0 8.568 0.024 8.928 ;
			RECT 0.0 8.952 0.024 9.312 ;
			RECT 0.0 9.336 0.024 9.696 ;
			RECT 0.0 9.72 0.024 10.08 ;
			RECT 0.0 10.104 0.024 10.464 ;
			RECT 0.0 10.488 0.024 10.848 ;
			RECT 0.0 10.872 0.024 11.232 ;
			RECT 0.0 11.256 0.024 11.616 ;
			RECT 0.0 11.64 0.024 11.664 ;
			RECT 0.0 11.688 0.024 12.048 ;
			RECT 0.0 12.072 0.024 12.432 ;
			RECT 0.0 12.456 0.024 12.816 ;
			RECT 0.0 12.84 0.024 13.2 ;
			RECT 0.0 13.224 0.024 13.584 ;
			RECT 0.0 13.608 0.024 13.968 ;
			RECT 0.0 13.992 0.024 14.352 ;
			RECT 0.0 14.376 0.024 14.736 ;
			RECT 0.0 14.76 0.024 15.12 ;
			RECT 0.0 15.144 0.024 15.504 ;
			RECT 0.0 15.528 0.024 15.888 ;
			RECT 0.0 15.912 0.024 16.272 ;
			RECT 0.0 16.296 0.024 16.656 ;
			RECT 0.0 16.68 0.024 17.04 ;
			RECT 0.0 17.064 0.024 17.424 ;
			RECT 0.0 17.448 0.024 17.472 ;
			RECT 0.0 17.496 0.024 17.856 ;
			RECT 0.0 17.88 0.024 18.24 ;
			RECT 0.0 18.264 0.024 18.624 ;
			RECT 0.0 18.648 0.024 19.008 ;
			RECT 0.0 19.032 0.024 19.392 ;
			RECT 0.0 19.416 0.024 19.776 ;
			RECT 0.0 19.8 0.024 20.16 ;
			RECT 0.0 20.184 0.024 20.208 ;
			RECT 0.0 20.232 0.024 20.592 ;
			RECT 0.0 20.616 0.024 20.976 ;
			RECT 0.0 16.8 0.024 21.0 ;

	END

END sram_asap7_16x256_1rw

MACRO sram_asap7_32x256_1rw
	CLASS BLOCK ;
	FOREIGN sram_asap7_32x256_1rw 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 16.72 BY 16.8 ;
	SYMMETRY X Y ;
	PIN clk
		DIRECTION INPUT ;
		USE CLOCK ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.408 0.024 15.432 ;

		END 

	END clk
	PIN rd_out[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.0 0.024 6.024 ;

		END 

	END rd_out[31]
	PIN rd_out[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.808 0.024 5.832 ;

		END 

	END rd_out[30]
	PIN rd_out[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.616 0.024 5.64 ;

		END 

	END rd_out[29]
	PIN rd_out[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.424 0.024 5.448 ;

		END 

	END rd_out[28]
	PIN rd_out[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.232 0.024 5.256 ;

		END 

	END rd_out[27]
	PIN rd_out[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.04 0.024 5.064 ;

		END 

	END rd_out[26]
	PIN rd_out[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.848 0.024 4.872 ;

		END 

	END rd_out[25]
	PIN rd_out[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.656 0.024 4.68 ;

		END 

	END rd_out[24]
	PIN rd_out[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.464 0.024 4.488 ;

		END 

	END rd_out[23]
	PIN rd_out[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.272 0.024 4.296 ;

		END 

	END rd_out[22]
	PIN rd_out[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.08 0.024 4.104 ;

		END 

	END rd_out[21]
	PIN rd_out[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.888 0.024 3.912 ;

		END 

	END rd_out[20]
	PIN rd_out[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.696 0.024 3.72 ;

		END 

	END rd_out[19]
	PIN rd_out[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.504 0.024 3.528 ;

		END 

	END rd_out[18]
	PIN rd_out[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.312 0.024 3.336 ;

		END 

	END rd_out[17]
	PIN rd_out[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.12 0.024 3.144 ;

		END 

	END rd_out[16]
	PIN rd_out[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.928 0.024 2.952 ;

		END 

	END rd_out[15]
	PIN rd_out[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.736 0.024 2.76 ;

		END 

	END rd_out[14]
	PIN rd_out[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.544 0.024 2.568 ;

		END 

	END rd_out[13]
	PIN rd_out[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.352 0.024 2.376 ;

		END 

	END rd_out[12]
	PIN rd_out[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.16 0.024 2.184 ;

		END 

	END rd_out[11]
	PIN rd_out[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.968 0.024 1.992 ;

		END 

	END rd_out[10]
	PIN rd_out[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.776 0.024 1.8 ;

		END 

	END rd_out[9]
	PIN rd_out[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.584 0.024 1.608 ;

		END 

	END rd_out[8]
	PIN rd_out[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.392 0.024 1.416 ;

		END 

	END rd_out[7]
	PIN rd_out[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.2 0.024 1.224 ;

		END 

	END rd_out[6]
	PIN rd_out[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.008 0.024 1.032 ;

		END 

	END rd_out[5]
	PIN rd_out[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.816 0.024 0.84 ;

		END 

	END rd_out[4]
	PIN rd_out[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.624 0.024 0.648 ;

		END 

	END rd_out[3]
	PIN rd_out[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.432 0.024 0.456 ;

		END 

	END rd_out[2]
	PIN rd_out[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.24 0.024 0.264 ;

		END 

	END rd_out[1]
	PIN rd_out[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.048 0.024 0.072 ;

		END 

	END rd_out[0]
	PIN we_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.024 0.024 15.048 ;

		END 

	END we_in
	PIN ce_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.216 0.024 15.24 ;

		END 

	END ce_in
	PIN addr_in[7]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.448 0.024 14.472 ;

		END 

	END addr_in[7]
	PIN addr_in[6]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.256 0.024 14.28 ;

		END 

	END addr_in[6]
	PIN addr_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.064 0.024 14.088 ;

		END 

	END addr_in[5]
	PIN addr_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.872 0.024 13.896 ;

		END 

	END addr_in[4]
	PIN addr_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.68 0.024 13.704 ;

		END 

	END addr_in[3]
	PIN addr_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.488 0.024 13.512 ;

		END 

	END addr_in[2]
	PIN addr_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.296 0.024 13.32 ;

		END 

	END addr_in[1]
	PIN addr_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.104 0.024 13.128 ;

		END 

	END addr_in[0]
	PIN wd_in[31]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.528 0.024 12.552 ;

		END 

	END wd_in[31]
	PIN wd_in[30]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.336 0.024 12.36 ;

		END 

	END wd_in[30]
	PIN wd_in[29]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.144 0.024 12.168 ;

		END 

	END wd_in[29]
	PIN wd_in[28]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.952 0.024 11.976 ;

		END 

	END wd_in[28]
	PIN wd_in[27]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.76 0.024 11.784 ;

		END 

	END wd_in[27]
	PIN wd_in[26]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.568 0.024 11.592 ;

		END 

	END wd_in[26]
	PIN wd_in[25]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.376 0.024 11.4 ;

		END 

	END wd_in[25]
	PIN wd_in[24]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.184 0.024 11.208 ;

		END 

	END wd_in[24]
	PIN wd_in[23]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.992 0.024 11.016 ;

		END 

	END wd_in[23]
	PIN wd_in[22]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.8 0.024 10.824 ;

		END 

	END wd_in[22]
	PIN wd_in[21]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.608 0.024 10.632 ;

		END 

	END wd_in[21]
	PIN wd_in[20]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.416 0.024 10.44 ;

		END 

	END wd_in[20]
	PIN wd_in[19]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.224 0.024 10.248 ;

		END 

	END wd_in[19]
	PIN wd_in[18]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.032 0.024 10.056 ;

		END 

	END wd_in[18]
	PIN wd_in[17]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.84 0.024 9.864 ;

		END 

	END wd_in[17]
	PIN wd_in[16]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.648 0.024 9.672 ;

		END 

	END wd_in[16]
	PIN wd_in[15]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.456 0.024 9.48 ;

		END 

	END wd_in[15]
	PIN wd_in[14]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.264 0.024 9.288 ;

		END 

	END wd_in[14]
	PIN wd_in[13]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.072 0.024 9.096 ;

		END 

	END wd_in[13]
	PIN wd_in[12]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.88 0.024 8.904 ;

		END 

	END wd_in[12]
	PIN wd_in[11]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.688 0.024 8.712 ;

		END 

	END wd_in[11]
	PIN wd_in[10]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.496 0.024 8.52 ;

		END 

	END wd_in[10]
	PIN wd_in[9]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.304 0.024 8.328 ;

		END 

	END wd_in[9]
	PIN wd_in[8]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.112 0.024 8.136 ;

		END 

	END wd_in[8]
	PIN wd_in[7]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.92 0.024 7.944 ;

		END 

	END wd_in[7]
	PIN wd_in[6]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.728 0.024 7.752 ;

		END 

	END wd_in[6]
	PIN wd_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.536 0.024 7.56 ;

		END 

	END wd_in[5]
	PIN wd_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.344 0.024 7.368 ;

		END 

	END wd_in[4]
	PIN wd_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.152 0.024 7.176 ;

		END 

	END wd_in[3]
	PIN wd_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.96 0.024 6.984 ;

		END 

	END wd_in[2]
	PIN wd_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.768 0.024 6.792 ;

		END 

	END wd_in[1]
	PIN wd_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.576 0.024 6.6 ;

		END 

	END wd_in[0]
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.0 16.672 0.096 ;
			RECT 0.048 0.768 16.672 0.864 ;
			RECT 0.048 1.536 16.672 1.632 ;
			RECT 0.048 2.304 16.672 2.4 ;
			RECT 0.048 3.072 16.672 3.168 ;
			RECT 0.048 3.84 16.672 3.936 ;
			RECT 0.048 4.608 16.672 4.704 ;
			RECT 0.048 5.376 16.672 5.472 ;
			RECT 0.048 6.144 16.672 6.24 ;
			RECT 0.048 6.912 16.672 7.008 ;
			RECT 0.048 7.68 16.672 7.776 ;
			RECT 0.048 8.448 16.672 8.544 ;
			RECT 0.048 9.216 16.672 9.312 ;
			RECT 0.048 9.984 16.672 10.08 ;
			RECT 0.048 10.752 16.672 10.848 ;
			RECT 0.048 11.52 16.672 11.616 ;
			RECT 0.048 12.288 16.672 12.384 ;
			RECT 0.048 13.056 16.672 13.152 ;
			RECT 0.048 13.824 16.672 13.92 ;
			RECT 0.048 14.592 16.672 14.688 ;
			RECT 0.048 15.36 16.672 15.456 ;
			RECT 0.048 16.128 16.672 16.224 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.384 16.672 0.48 ;
			RECT 0.048 1.152 16.672 1.248 ;
			RECT 0.048 1.92 16.672 2.016 ;
			RECT 0.048 2.688 16.672 2.784 ;
			RECT 0.048 3.456 16.672 3.552 ;
			RECT 0.048 4.224 16.672 4.32 ;
			RECT 0.048 4.992 16.672 5.088 ;
			RECT 0.048 5.76 16.672 5.856 ;
			RECT 0.048 6.528 16.672 6.624 ;
			RECT 0.048 7.296 16.672 7.392 ;
			RECT 0.048 8.064 16.672 8.16 ;
			RECT 0.048 8.832 16.672 8.928 ;
			RECT 0.048 9.6 16.672 9.696 ;
			RECT 0.048 10.368 16.672 10.464 ;
			RECT 0.048 11.136 16.672 11.232 ;
			RECT 0.048 11.904 16.672 12.0 ;
			RECT 0.048 12.672 16.672 12.768 ;
			RECT 0.048 13.44 16.672 13.536 ;
			RECT 0.048 14.208 16.672 14.304 ;
			RECT 0.048 14.976 16.672 15.072 ;
			RECT 0.048 15.744 16.672 15.84 ;
			RECT 0.048 16.512 16.672 16.608 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.0 0.0 16.72 16.8 ;
			LAYER M2 ;
			RECT 0.0 0.0 16.72 16.8 ;
			LAYER M3 ;
			RECT 0.0 0.0 16.72 16.8 ;
			LAYER M4 ;
			RECT 0.024 0.0 0.048 16.8 ;
			RECT 16.672 0.0 16.72 16.8 ;
			RECT 0.048 0.0 16.672 0.0 ;
			RECT 0.048 0.096 16.672 0.384 ;
			RECT 0.048 0.48 16.672 0.768 ;
			RECT 0.048 0.864 16.672 1.152 ;
			RECT 0.048 1.248 16.672 1.536 ;
			RECT 0.048 1.632 16.672 1.92 ;
			RECT 0.048 2.016 16.672 2.304 ;
			RECT 0.048 2.4 16.672 2.688 ;
			RECT 0.048 2.784 16.672 3.072 ;
			RECT 0.048 3.168 16.672 3.456 ;
			RECT 0.048 3.552 16.672 3.84 ;
			RECT 0.048 3.936 16.672 4.224 ;
			RECT 0.048 4.32 16.672 4.608 ;
			RECT 0.048 4.704 16.672 4.992 ;
			RECT 0.048 5.088 16.672 5.376 ;
			RECT 0.048 5.472 16.672 5.76 ;
			RECT 0.048 5.856 16.672 6.144 ;
			RECT 0.048 6.24 16.672 6.528 ;
			RECT 0.048 6.624 16.672 6.912 ;
			RECT 0.048 7.008 16.672 7.296 ;
			RECT 0.048 7.392 16.672 7.68 ;
			RECT 0.048 7.776 16.672 8.064 ;
			RECT 0.048 8.16 16.672 8.448 ;
			RECT 0.048 8.544 16.672 8.832 ;
			RECT 0.048 8.928 16.672 9.216 ;
			RECT 0.048 9.312 16.672 9.6 ;
			RECT 0.048 9.696 16.672 9.984 ;
			RECT 0.048 10.08 16.672 10.368 ;
			RECT 0.048 10.464 16.672 10.752 ;
			RECT 0.048 10.848 16.672 11.136 ;
			RECT 0.048 11.232 16.672 11.52 ;
			RECT 0.048 11.616 16.672 11.904 ;
			RECT 0.048 12.0 16.672 12.288 ;
			RECT 0.048 12.384 16.672 12.672 ;
			RECT 0.048 12.768 16.672 13.056 ;
			RECT 0.048 13.152 16.672 13.44 ;
			RECT 0.048 13.536 16.672 13.824 ;
			RECT 0.048 13.92 16.672 14.208 ;
			RECT 0.048 14.304 16.672 14.592 ;
			RECT 0.048 14.688 16.672 14.976 ;
			RECT 0.048 15.072 16.672 15.36 ;
			RECT 0.048 15.456 16.672 15.744 ;
			RECT 0.048 15.84 16.672 16.128 ;
			RECT 0.048 16.224 16.672 16.512 ;
			RECT 0.048 16.608 16.672 16.8 ;
			RECT 0.0 0.0 0.024 0.048 ;
			RECT 0.0 0.072 0.024 0.24 ;
			RECT 0.0 0.264 0.024 0.432 ;
			RECT 0.0 0.456 0.024 0.624 ;
			RECT 0.0 0.648 0.024 0.816 ;
			RECT 0.0 0.84 0.024 1.008 ;
			RECT 0.0 1.032 0.024 1.2 ;
			RECT 0.0 1.224 0.024 1.392 ;
			RECT 0.0 1.416 0.024 1.584 ;
			RECT 0.0 1.608 0.024 1.776 ;
			RECT 0.0 1.8 0.024 1.968 ;
			RECT 0.0 1.992 0.024 2.16 ;
			RECT 0.0 2.184 0.024 2.352 ;
			RECT 0.0 2.376 0.024 2.544 ;
			RECT 0.0 2.568 0.024 2.736 ;
			RECT 0.0 2.76 0.024 2.928 ;
			RECT 0.0 2.952 0.024 3.12 ;
			RECT 0.0 3.144 0.024 3.312 ;
			RECT 0.0 3.336 0.024 3.504 ;
			RECT 0.0 3.528 0.024 3.696 ;
			RECT 0.0 3.72 0.024 3.888 ;
			RECT 0.0 3.912 0.024 4.08 ;
			RECT 0.0 4.104 0.024 4.272 ;
			RECT 0.0 4.296 0.024 4.464 ;
			RECT 0.0 4.488 0.024 4.656 ;
			RECT 0.0 4.68 0.024 4.848 ;
			RECT 0.0 4.872 0.024 5.04 ;
			RECT 0.0 5.064 0.024 5.232 ;
			RECT 0.0 5.256 0.024 5.424 ;
			RECT 0.0 5.448 0.024 5.616 ;
			RECT 0.0 5.64 0.024 5.808 ;
			RECT 0.0 5.832 0.024 6.0 ;
			RECT 0.0 6.024 0.024 6.576 ;
			RECT 0.0 6.6 0.024 6.768 ;
			RECT 0.0 6.792 0.024 6.96 ;
			RECT 0.0 6.984 0.024 7.152 ;
			RECT 0.0 7.176 0.024 7.344 ;
			RECT 0.0 7.368 0.024 7.536 ;
			RECT 0.0 7.56 0.024 7.728 ;
			RECT 0.0 7.752 0.024 7.92 ;
			RECT 0.0 7.944 0.024 8.112 ;
			RECT 0.0 8.136 0.024 8.304 ;
			RECT 0.0 8.328 0.024 8.496 ;
			RECT 0.0 8.52 0.024 8.688 ;
			RECT 0.0 8.712 0.024 8.88 ;
			RECT 0.0 8.904 0.024 9.072 ;
			RECT 0.0 9.096 0.024 9.264 ;
			RECT 0.0 9.288 0.024 9.456 ;
			RECT 0.0 9.48 0.024 9.648 ;
			RECT 0.0 9.672 0.024 9.84 ;
			RECT 0.0 9.864 0.024 10.032 ;
			RECT 0.0 10.056 0.024 10.224 ;
			RECT 0.0 10.248 0.024 10.416 ;
			RECT 0.0 10.44 0.024 10.608 ;
			RECT 0.0 10.632 0.024 10.8 ;
			RECT 0.0 10.824 0.024 10.992 ;
			RECT 0.0 11.016 0.024 11.184 ;
			RECT 0.0 11.208 0.024 11.376 ;
			RECT 0.0 11.4 0.024 11.568 ;
			RECT 0.0 11.592 0.024 11.76 ;
			RECT 0.0 11.784 0.024 11.952 ;
			RECT 0.0 11.976 0.024 12.144 ;
			RECT 0.0 12.168 0.024 12.336 ;
			RECT 0.0 12.36 0.024 12.528 ;
			RECT 0.0 12.552 0.024 13.104 ;
			RECT 0.0 13.128 0.024 13.296 ;
			RECT 0.0 13.32 0.024 13.488 ;
			RECT 0.0 13.512 0.024 13.68 ;
			RECT 0.0 13.704 0.024 13.872 ;
			RECT 0.0 13.896 0.024 14.064 ;
			RECT 0.0 14.088 0.024 14.256 ;
			RECT 0.0 14.28 0.024 14.448 ;
			RECT 0.0 14.472 0.024 14.64 ;
			RECT 0.0 14.664 0.024 14.832 ;
			RECT 0.0 14.856 0.024 15.024 ;
			RECT 0.0 15.048 0.024 15.216 ;
			RECT 0.0 15.24 0.024 15.408 ;
			RECT 0.0 15.432 0.024 15.6 ;
			RECT 0.0 15.624 0.024 15.792 ;
			RECT 0.0 15.816 0.024 15.984 ;
			RECT 0.0 16.008 0.024 16.176 ;
			RECT 0.0 16.2 0.024 16.368 ;
			RECT 0.0 16.392 0.024 16.56 ;
			RECT 0.0 16.584 0.024 16.752 ;
			RECT 0.0 16.776 0.024 16.944 ;
			RECT 0.0 16.968 0.024 17.136 ;
			RECT 0.0 17.16 0.024 17.328 ;
			RECT 0.0 17.352 0.024 17.52 ;
			RECT 0.0 17.544 0.024 17.712 ;
			RECT 0.0 17.736 0.024 17.904 ;
			RECT 0.0 17.928 0.024 18.096 ;
			RECT 0.0 18.12 0.024 18.288 ;
			RECT 0.0 18.312 0.024 18.48 ;
			RECT 0.0 18.504 0.024 18.672 ;
			RECT 0.0 18.696 0.024 18.864 ;
			RECT 0.0 18.888 0.024 19.056 ;
			RECT 0.0 19.08 0.024 19.632 ;
			RECT 0.0 19.656 0.024 19.824 ;
			RECT 0.0 19.848 0.024 20.016 ;
			RECT 0.0 20.04 0.024 20.208 ;
			RECT 0.0 20.232 0.024 20.4 ;
			RECT 0.0 20.424 0.024 20.592 ;
			RECT 0.0 20.616 0.024 20.784 ;
			RECT 0.0 20.808 0.024 20.976 ;
			RECT 0.0 21.0 0.024 21.552 ;
			RECT 0.0 21.576 0.024 21.744 ;
			RECT 0.0 21.768 0.024 21.936 ;
			RECT 0.0 16.8 0.024 21.96 ;

	END

END sram_asap7_32x256_1rw

MACRO sram_asap7_64x256_1rw
	CLASS BLOCK ;
	FOREIGN sram_asap7_64x256_1rw 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 16.72 BY 33.6 ;
	SYMMETRY X Y ;
	PIN clk
		DIRECTION INPUT ;
		USE CLOCK ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 32.592 0.024 32.616 ;

		END 

	END clk
	PIN rd_out[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.168 0.024 15.192 ;

		END 

	END rd_out[63]
	PIN rd_out[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.928 0.024 14.952 ;

		END 

	END rd_out[62]
	PIN rd_out[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.688 0.024 14.712 ;

		END 

	END rd_out[61]
	PIN rd_out[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.448 0.024 14.472 ;

		END 

	END rd_out[60]
	PIN rd_out[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.208 0.024 14.232 ;

		END 

	END rd_out[59]
	PIN rd_out[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.968 0.024 13.992 ;

		END 

	END rd_out[58]
	PIN rd_out[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.728 0.024 13.752 ;

		END 

	END rd_out[57]
	PIN rd_out[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.488 0.024 13.512 ;

		END 

	END rd_out[56]
	PIN rd_out[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.248 0.024 13.272 ;

		END 

	END rd_out[55]
	PIN rd_out[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.008 0.024 13.032 ;

		END 

	END rd_out[54]
	PIN rd_out[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.768 0.024 12.792 ;

		END 

	END rd_out[53]
	PIN rd_out[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.528 0.024 12.552 ;

		END 

	END rd_out[52]
	PIN rd_out[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.288 0.024 12.312 ;

		END 

	END rd_out[51]
	PIN rd_out[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.048 0.024 12.072 ;

		END 

	END rd_out[50]
	PIN rd_out[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.808 0.024 11.832 ;

		END 

	END rd_out[49]
	PIN rd_out[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.568 0.024 11.592 ;

		END 

	END rd_out[48]
	PIN rd_out[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.328 0.024 11.352 ;

		END 

	END rd_out[47]
	PIN rd_out[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.088 0.024 11.112 ;

		END 

	END rd_out[46]
	PIN rd_out[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.848 0.024 10.872 ;

		END 

	END rd_out[45]
	PIN rd_out[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.608 0.024 10.632 ;

		END 

	END rd_out[44]
	PIN rd_out[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.368 0.024 10.392 ;

		END 

	END rd_out[43]
	PIN rd_out[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.128 0.024 10.152 ;

		END 

	END rd_out[42]
	PIN rd_out[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.888 0.024 9.912 ;

		END 

	END rd_out[41]
	PIN rd_out[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.648 0.024 9.672 ;

		END 

	END rd_out[40]
	PIN rd_out[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.408 0.024 9.432 ;

		END 

	END rd_out[39]
	PIN rd_out[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.168 0.024 9.192 ;

		END 

	END rd_out[38]
	PIN rd_out[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.928 0.024 8.952 ;

		END 

	END rd_out[37]
	PIN rd_out[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.688 0.024 8.712 ;

		END 

	END rd_out[36]
	PIN rd_out[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.448 0.024 8.472 ;

		END 

	END rd_out[35]
	PIN rd_out[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.208 0.024 8.232 ;

		END 

	END rd_out[34]
	PIN rd_out[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.968 0.024 7.992 ;

		END 

	END rd_out[33]
	PIN rd_out[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.728 0.024 7.752 ;

		END 

	END rd_out[32]
	PIN rd_out[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.488 0.024 7.512 ;

		END 

	END rd_out[31]
	PIN rd_out[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.248 0.024 7.272 ;

		END 

	END rd_out[30]
	PIN rd_out[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.008 0.024 7.032 ;

		END 

	END rd_out[29]
	PIN rd_out[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.768 0.024 6.792 ;

		END 

	END rd_out[28]
	PIN rd_out[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.528 0.024 6.552 ;

		END 

	END rd_out[27]
	PIN rd_out[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.288 0.024 6.312 ;

		END 

	END rd_out[26]
	PIN rd_out[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.048 0.024 6.072 ;

		END 

	END rd_out[25]
	PIN rd_out[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.808 0.024 5.832 ;

		END 

	END rd_out[24]
	PIN rd_out[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.568 0.024 5.592 ;

		END 

	END rd_out[23]
	PIN rd_out[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.328 0.024 5.352 ;

		END 

	END rd_out[22]
	PIN rd_out[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.088 0.024 5.112 ;

		END 

	END rd_out[21]
	PIN rd_out[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.848 0.024 4.872 ;

		END 

	END rd_out[20]
	PIN rd_out[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.608 0.024 4.632 ;

		END 

	END rd_out[19]
	PIN rd_out[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.368 0.024 4.392 ;

		END 

	END rd_out[18]
	PIN rd_out[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.128 0.024 4.152 ;

		END 

	END rd_out[17]
	PIN rd_out[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.888 0.024 3.912 ;

		END 

	END rd_out[16]
	PIN rd_out[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.648 0.024 3.672 ;

		END 

	END rd_out[15]
	PIN rd_out[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.408 0.024 3.432 ;

		END 

	END rd_out[14]
	PIN rd_out[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.168 0.024 3.192 ;

		END 

	END rd_out[13]
	PIN rd_out[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.928 0.024 2.952 ;

		END 

	END rd_out[12]
	PIN rd_out[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.688 0.024 2.712 ;

		END 

	END rd_out[11]
	PIN rd_out[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.448 0.024 2.472 ;

		END 

	END rd_out[10]
	PIN rd_out[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.208 0.024 2.232 ;

		END 

	END rd_out[9]
	PIN rd_out[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.968 0.024 1.992 ;

		END 

	END rd_out[8]
	PIN rd_out[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.728 0.024 1.752 ;

		END 

	END rd_out[7]
	PIN rd_out[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.488 0.024 1.512 ;

		END 

	END rd_out[6]
	PIN rd_out[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.248 0.024 1.272 ;

		END 

	END rd_out[5]
	PIN rd_out[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.008 0.024 1.032 ;

		END 

	END rd_out[4]
	PIN rd_out[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.768 0.024 0.792 ;

		END 

	END rd_out[3]
	PIN rd_out[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.528 0.024 0.552 ;

		END 

	END rd_out[2]
	PIN rd_out[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.288 0.024 0.312 ;

		END 

	END rd_out[1]
	PIN rd_out[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.048 0.024 0.072 ;

		END 

	END rd_out[0]
	PIN we_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 32.112 0.024 32.136 ;

		END 

	END we_in
	PIN ce_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 32.352 0.024 32.376 ;

		END 

	END ce_in
	PIN addr_in[7]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 32.064 0.024 32.088 ;

		END 

	END addr_in[7]
	PIN addr_in[6]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 31.824 0.024 31.848 ;

		END 

	END addr_in[6]
	PIN addr_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 31.584 0.024 31.608 ;

		END 

	END addr_in[5]
	PIN addr_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 31.344 0.024 31.368 ;

		END 

	END addr_in[4]
	PIN addr_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 31.104 0.024 31.128 ;

		END 

	END addr_in[3]
	PIN addr_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 30.864 0.024 30.888 ;

		END 

	END addr_in[2]
	PIN addr_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 30.624 0.024 30.648 ;

		END 

	END addr_in[1]
	PIN addr_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 30.384 0.024 30.408 ;

		END 

	END addr_in[0]
	PIN wd_in[63]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 30.336 0.024 30.36 ;

		END 

	END wd_in[63]
	PIN wd_in[62]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 30.096 0.024 30.12 ;

		END 

	END wd_in[62]
	PIN wd_in[61]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 29.856 0.024 29.88 ;

		END 

	END wd_in[61]
	PIN wd_in[60]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 29.616 0.024 29.64 ;

		END 

	END wd_in[60]
	PIN wd_in[59]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 29.376 0.024 29.4 ;

		END 

	END wd_in[59]
	PIN wd_in[58]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 29.136 0.024 29.16 ;

		END 

	END wd_in[58]
	PIN wd_in[57]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 28.896 0.024 28.92 ;

		END 

	END wd_in[57]
	PIN wd_in[56]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 28.656 0.024 28.68 ;

		END 

	END wd_in[56]
	PIN wd_in[55]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 28.416 0.024 28.44 ;

		END 

	END wd_in[55]
	PIN wd_in[54]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 28.176 0.024 28.2 ;

		END 

	END wd_in[54]
	PIN wd_in[53]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 27.936 0.024 27.96 ;

		END 

	END wd_in[53]
	PIN wd_in[52]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 27.696 0.024 27.72 ;

		END 

	END wd_in[52]
	PIN wd_in[51]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 27.456 0.024 27.48 ;

		END 

	END wd_in[51]
	PIN wd_in[50]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 27.216 0.024 27.24 ;

		END 

	END wd_in[50]
	PIN wd_in[49]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 26.976 0.024 27.0 ;

		END 

	END wd_in[49]
	PIN wd_in[48]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 26.736 0.024 26.76 ;

		END 

	END wd_in[48]
	PIN wd_in[47]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 26.496 0.024 26.52 ;

		END 

	END wd_in[47]
	PIN wd_in[46]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 26.256 0.024 26.28 ;

		END 

	END wd_in[46]
	PIN wd_in[45]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 26.016 0.024 26.04 ;

		END 

	END wd_in[45]
	PIN wd_in[44]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 25.776 0.024 25.8 ;

		END 

	END wd_in[44]
	PIN wd_in[43]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 25.536 0.024 25.56 ;

		END 

	END wd_in[43]
	PIN wd_in[42]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 25.296 0.024 25.32 ;

		END 

	END wd_in[42]
	PIN wd_in[41]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 25.056 0.024 25.08 ;

		END 

	END wd_in[41]
	PIN wd_in[40]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 24.816 0.024 24.84 ;

		END 

	END wd_in[40]
	PIN wd_in[39]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 24.576 0.024 24.6 ;

		END 

	END wd_in[39]
	PIN wd_in[38]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 24.336 0.024 24.36 ;

		END 

	END wd_in[38]
	PIN wd_in[37]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 24.096 0.024 24.12 ;

		END 

	END wd_in[37]
	PIN wd_in[36]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 23.856 0.024 23.88 ;

		END 

	END wd_in[36]
	PIN wd_in[35]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 23.616 0.024 23.64 ;

		END 

	END wd_in[35]
	PIN wd_in[34]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 23.376 0.024 23.4 ;

		END 

	END wd_in[34]
	PIN wd_in[33]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 23.136 0.024 23.16 ;

		END 

	END wd_in[33]
	PIN wd_in[32]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 22.896 0.024 22.92 ;

		END 

	END wd_in[32]
	PIN wd_in[31]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 22.656 0.024 22.68 ;

		END 

	END wd_in[31]
	PIN wd_in[30]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 22.416 0.024 22.44 ;

		END 

	END wd_in[30]
	PIN wd_in[29]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 22.176 0.024 22.2 ;

		END 

	END wd_in[29]
	PIN wd_in[28]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 21.936 0.024 21.96 ;

		END 

	END wd_in[28]
	PIN wd_in[27]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 21.696 0.024 21.72 ;

		END 

	END wd_in[27]
	PIN wd_in[26]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 21.456 0.024 21.48 ;

		END 

	END wd_in[26]
	PIN wd_in[25]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 21.216 0.024 21.24 ;

		END 

	END wd_in[25]
	PIN wd_in[24]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 20.976 0.024 21.0 ;

		END 

	END wd_in[24]
	PIN wd_in[23]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 20.736 0.024 20.76 ;

		END 

	END wd_in[23]
	PIN wd_in[22]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 20.496 0.024 20.52 ;

		END 

	END wd_in[22]
	PIN wd_in[21]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 20.256 0.024 20.28 ;

		END 

	END wd_in[21]
	PIN wd_in[20]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 20.016 0.024 20.04 ;

		END 

	END wd_in[20]
	PIN wd_in[19]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 19.776 0.024 19.8 ;

		END 

	END wd_in[19]
	PIN wd_in[18]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 19.536 0.024 19.56 ;

		END 

	END wd_in[18]
	PIN wd_in[17]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 19.296 0.024 19.32 ;

		END 

	END wd_in[17]
	PIN wd_in[16]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 19.056 0.024 19.08 ;

		END 

	END wd_in[16]
	PIN wd_in[15]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 18.816 0.024 18.84 ;

		END 

	END wd_in[15]
	PIN wd_in[14]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 18.576 0.024 18.6 ;

		END 

	END wd_in[14]
	PIN wd_in[13]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 18.336 0.024 18.36 ;

		END 

	END wd_in[13]
	PIN wd_in[12]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 18.096 0.024 18.12 ;

		END 

	END wd_in[12]
	PIN wd_in[11]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 17.856 0.024 17.88 ;

		END 

	END wd_in[11]
	PIN wd_in[10]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 17.616 0.024 17.64 ;

		END 

	END wd_in[10]
	PIN wd_in[9]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 17.376 0.024 17.4 ;

		END 

	END wd_in[9]
	PIN wd_in[8]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 17.136 0.024 17.16 ;

		END 

	END wd_in[8]
	PIN wd_in[7]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 16.896 0.024 16.92 ;

		END 

	END wd_in[7]
	PIN wd_in[6]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 16.656 0.024 16.68 ;

		END 

	END wd_in[6]
	PIN wd_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 16.416 0.024 16.44 ;

		END 

	END wd_in[5]
	PIN wd_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 16.176 0.024 16.2 ;

		END 

	END wd_in[4]
	PIN wd_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.936 0.024 15.96 ;

		END 

	END wd_in[3]
	PIN wd_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.696 0.024 15.72 ;

		END 

	END wd_in[2]
	PIN wd_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.456 0.024 15.48 ;

		END 

	END wd_in[1]
	PIN wd_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.216 0.024 15.24 ;

		END 

	END wd_in[0]
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.0 16.672 0.096 ;
			RECT 0.048 0.768 16.672 0.864 ;
			RECT 0.048 1.536 16.672 1.632 ;
			RECT 0.048 2.304 16.672 2.4 ;
			RECT 0.048 3.072 16.672 3.168 ;
			RECT 0.048 3.84 16.672 3.936 ;
			RECT 0.048 4.608 16.672 4.704 ;
			RECT 0.048 5.376 16.672 5.472 ;
			RECT 0.048 6.144 16.672 6.24 ;
			RECT 0.048 6.912 16.672 7.008 ;
			RECT 0.048 7.68 16.672 7.776 ;
			RECT 0.048 8.448 16.672 8.544 ;
			RECT 0.048 9.216 16.672 9.312 ;
			RECT 0.048 9.984 16.672 10.08 ;
			RECT 0.048 10.752 16.672 10.848 ;
			RECT 0.048 11.52 16.672 11.616 ;
			RECT 0.048 12.288 16.672 12.384 ;
			RECT 0.048 13.056 16.672 13.152 ;
			RECT 0.048 13.824 16.672 13.92 ;
			RECT 0.048 14.592 16.672 14.688 ;
			RECT 0.048 15.36 16.672 15.456 ;
			RECT 0.048 16.128 16.672 16.224 ;
			RECT 0.048 16.896 16.672 16.992 ;
			RECT 0.048 17.664 16.672 17.76 ;
			RECT 0.048 18.432 16.672 18.528 ;
			RECT 0.048 19.2 16.672 19.296 ;
			RECT 0.048 19.968 16.672 20.064 ;
			RECT 0.048 20.736 16.672 20.832 ;
			RECT 0.048 21.504 16.672 21.6 ;
			RECT 0.048 22.272 16.672 22.368 ;
			RECT 0.048 23.04 16.672 23.136 ;
			RECT 0.048 23.808 16.672 23.904 ;
			RECT 0.048 24.576 16.672 24.672 ;
			RECT 0.048 25.344 16.672 25.44 ;
			RECT 0.048 26.112 16.672 26.208 ;
			RECT 0.048 26.88 16.672 26.976 ;
			RECT 0.048 27.648 16.672 27.744 ;
			RECT 0.048 28.416 16.672 28.512 ;
			RECT 0.048 29.184 16.672 29.28 ;
			RECT 0.048 29.952 16.672 30.048 ;
			RECT 0.048 30.72 16.672 30.816 ;
			RECT 0.048 31.488 16.672 31.584 ;
			RECT 0.048 32.256 16.672 32.352 ;
			RECT 0.048 33.024 16.672 33.12 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.384 16.672 0.48 ;
			RECT 0.048 1.152 16.672 1.248 ;
			RECT 0.048 1.92 16.672 2.016 ;
			RECT 0.048 2.688 16.672 2.784 ;
			RECT 0.048 3.456 16.672 3.552 ;
			RECT 0.048 4.224 16.672 4.32 ;
			RECT 0.048 4.992 16.672 5.088 ;
			RECT 0.048 5.76 16.672 5.856 ;
			RECT 0.048 6.528 16.672 6.624 ;
			RECT 0.048 7.296 16.672 7.392 ;
			RECT 0.048 8.064 16.672 8.16 ;
			RECT 0.048 8.832 16.672 8.928 ;
			RECT 0.048 9.6 16.672 9.696 ;
			RECT 0.048 10.368 16.672 10.464 ;
			RECT 0.048 11.136 16.672 11.232 ;
			RECT 0.048 11.904 16.672 12.0 ;
			RECT 0.048 12.672 16.672 12.768 ;
			RECT 0.048 13.44 16.672 13.536 ;
			RECT 0.048 14.208 16.672 14.304 ;
			RECT 0.048 14.976 16.672 15.072 ;
			RECT 0.048 15.744 16.672 15.84 ;
			RECT 0.048 16.512 16.672 16.608 ;
			RECT 0.048 17.28 16.672 17.376 ;
			RECT 0.048 18.048 16.672 18.144 ;
			RECT 0.048 18.816 16.672 18.912 ;
			RECT 0.048 19.584 16.672 19.68 ;
			RECT 0.048 20.352 16.672 20.448 ;
			RECT 0.048 21.12 16.672 21.216 ;
			RECT 0.048 21.888 16.672 21.984 ;
			RECT 0.048 22.656 16.672 22.752 ;
			RECT 0.048 23.424 16.672 23.52 ;
			RECT 0.048 24.192 16.672 24.288 ;
			RECT 0.048 24.96 16.672 25.056 ;
			RECT 0.048 25.728 16.672 25.824 ;
			RECT 0.048 26.496 16.672 26.592 ;
			RECT 0.048 27.264 16.672 27.36 ;
			RECT 0.048 28.032 16.672 28.128 ;
			RECT 0.048 28.8 16.672 28.896 ;
			RECT 0.048 29.568 16.672 29.664 ;
			RECT 0.048 30.336 16.672 30.432 ;
			RECT 0.048 31.104 16.672 31.2 ;
			RECT 0.048 31.872 16.672 31.968 ;
			RECT 0.048 32.64 16.672 32.736 ;
			RECT 0.048 33.408 16.672 33.504 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.0 0.0 16.72 33.6 ;
			LAYER M2 ;
			RECT 0.0 0.0 16.72 33.6 ;
			LAYER M3 ;
			RECT 0.0 0.0 16.72 33.6 ;
			LAYER M4 ;
			RECT 0.024 0.0 0.048 33.6 ;
			RECT 16.672 0.0 16.72 33.6 ;
			RECT 0.048 0.0 16.672 0.0 ;
			RECT 0.048 0.096 16.672 0.384 ;
			RECT 0.048 0.48 16.672 0.768 ;
			RECT 0.048 0.864 16.672 1.152 ;
			RECT 0.048 1.248 16.672 1.536 ;
			RECT 0.048 1.632 16.672 1.92 ;
			RECT 0.048 2.016 16.672 2.304 ;
			RECT 0.048 2.4 16.672 2.688 ;
			RECT 0.048 2.784 16.672 3.072 ;
			RECT 0.048 3.168 16.672 3.456 ;
			RECT 0.048 3.552 16.672 3.84 ;
			RECT 0.048 3.936 16.672 4.224 ;
			RECT 0.048 4.32 16.672 4.608 ;
			RECT 0.048 4.704 16.672 4.992 ;
			RECT 0.048 5.088 16.672 5.376 ;
			RECT 0.048 5.472 16.672 5.76 ;
			RECT 0.048 5.856 16.672 6.144 ;
			RECT 0.048 6.24 16.672 6.528 ;
			RECT 0.048 6.624 16.672 6.912 ;
			RECT 0.048 7.008 16.672 7.296 ;
			RECT 0.048 7.392 16.672 7.68 ;
			RECT 0.048 7.776 16.672 8.064 ;
			RECT 0.048 8.16 16.672 8.448 ;
			RECT 0.048 8.544 16.672 8.832 ;
			RECT 0.048 8.928 16.672 9.216 ;
			RECT 0.048 9.312 16.672 9.6 ;
			RECT 0.048 9.696 16.672 9.984 ;
			RECT 0.048 10.08 16.672 10.368 ;
			RECT 0.048 10.464 16.672 10.752 ;
			RECT 0.048 10.848 16.672 11.136 ;
			RECT 0.048 11.232 16.672 11.52 ;
			RECT 0.048 11.616 16.672 11.904 ;
			RECT 0.048 12.0 16.672 12.288 ;
			RECT 0.048 12.384 16.672 12.672 ;
			RECT 0.048 12.768 16.672 13.056 ;
			RECT 0.048 13.152 16.672 13.44 ;
			RECT 0.048 13.536 16.672 13.824 ;
			RECT 0.048 13.92 16.672 14.208 ;
			RECT 0.048 14.304 16.672 14.592 ;
			RECT 0.048 14.688 16.672 14.976 ;
			RECT 0.048 15.072 16.672 15.36 ;
			RECT 0.048 15.456 16.672 15.744 ;
			RECT 0.048 15.84 16.672 16.128 ;
			RECT 0.048 16.224 16.672 16.512 ;
			RECT 0.048 16.608 16.672 16.896 ;
			RECT 0.048 16.992 16.672 17.28 ;
			RECT 0.048 17.376 16.672 17.664 ;
			RECT 0.048 17.76 16.672 18.048 ;
			RECT 0.048 18.144 16.672 18.432 ;
			RECT 0.048 18.528 16.672 18.816 ;
			RECT 0.048 18.912 16.672 19.2 ;
			RECT 0.048 19.296 16.672 19.584 ;
			RECT 0.048 19.68 16.672 19.968 ;
			RECT 0.048 20.064 16.672 20.352 ;
			RECT 0.048 20.448 16.672 20.736 ;
			RECT 0.048 20.832 16.672 21.12 ;
			RECT 0.048 21.216 16.672 21.504 ;
			RECT 0.048 21.6 16.672 21.888 ;
			RECT 0.048 21.984 16.672 22.272 ;
			RECT 0.048 22.368 16.672 22.656 ;
			RECT 0.048 22.752 16.672 23.04 ;
			RECT 0.048 23.136 16.672 23.424 ;
			RECT 0.048 23.52 16.672 23.808 ;
			RECT 0.048 23.904 16.672 24.192 ;
			RECT 0.048 24.288 16.672 24.576 ;
			RECT 0.048 24.672 16.672 24.96 ;
			RECT 0.048 25.056 16.672 25.344 ;
			RECT 0.048 25.44 16.672 25.728 ;
			RECT 0.048 25.824 16.672 26.112 ;
			RECT 0.048 26.208 16.672 26.496 ;
			RECT 0.048 26.592 16.672 26.88 ;
			RECT 0.048 26.976 16.672 27.264 ;
			RECT 0.048 27.36 16.672 27.648 ;
			RECT 0.048 27.744 16.672 28.032 ;
			RECT 0.048 28.128 16.672 28.416 ;
			RECT 0.048 28.512 16.672 28.8 ;
			RECT 0.048 28.896 16.672 29.184 ;
			RECT 0.048 29.28 16.672 29.568 ;
			RECT 0.048 29.664 16.672 29.952 ;
			RECT 0.048 30.048 16.672 30.336 ;
			RECT 0.048 30.432 16.672 30.72 ;
			RECT 0.048 30.816 16.672 31.104 ;
			RECT 0.048 31.2 16.672 31.488 ;
			RECT 0.048 31.584 16.672 31.872 ;
			RECT 0.048 31.968 16.672 32.256 ;
			RECT 0.048 32.352 16.672 32.64 ;
			RECT 0.048 32.736 16.672 33.024 ;
			RECT 0.048 33.12 16.672 33.408 ;
			RECT 0.048 33.504 16.672 33.6 ;
			RECT 0.0 0.0 0.024 0.048 ;
			RECT 0.0 0.072 0.024 0.288 ;
			RECT 0.0 0.312 0.024 0.528 ;
			RECT 0.0 0.552 0.024 0.768 ;
			RECT 0.0 0.792 0.024 1.008 ;
			RECT 0.0 1.032 0.024 1.248 ;
			RECT 0.0 1.272 0.024 1.488 ;
			RECT 0.0 1.512 0.024 1.728 ;
			RECT 0.0 1.752 0.024 1.968 ;
			RECT 0.0 1.992 0.024 2.208 ;
			RECT 0.0 2.232 0.024 2.448 ;
			RECT 0.0 2.472 0.024 2.688 ;
			RECT 0.0 2.712 0.024 2.928 ;
			RECT 0.0 2.952 0.024 3.168 ;
			RECT 0.0 3.192 0.024 3.408 ;
			RECT 0.0 3.432 0.024 3.648 ;
			RECT 0.0 3.672 0.024 3.888 ;
			RECT 0.0 3.912 0.024 4.128 ;
			RECT 0.0 4.152 0.024 4.368 ;
			RECT 0.0 4.392 0.024 4.608 ;
			RECT 0.0 4.632 0.024 4.848 ;
			RECT 0.0 4.872 0.024 5.088 ;
			RECT 0.0 5.112 0.024 5.328 ;
			RECT 0.0 5.352 0.024 5.568 ;
			RECT 0.0 5.592 0.024 5.808 ;
			RECT 0.0 5.832 0.024 6.048 ;
			RECT 0.0 6.072 0.024 6.288 ;
			RECT 0.0 6.312 0.024 6.528 ;
			RECT 0.0 6.552 0.024 6.768 ;
			RECT 0.0 6.792 0.024 7.008 ;
			RECT 0.0 7.032 0.024 7.248 ;
			RECT 0.0 7.272 0.024 7.488 ;
			RECT 0.0 7.512 0.024 7.728 ;
			RECT 0.0 7.752 0.024 7.968 ;
			RECT 0.0 7.992 0.024 8.208 ;
			RECT 0.0 8.232 0.024 8.448 ;
			RECT 0.0 8.472 0.024 8.688 ;
			RECT 0.0 8.712 0.024 8.928 ;
			RECT 0.0 8.952 0.024 9.168 ;
			RECT 0.0 9.192 0.024 9.408 ;
			RECT 0.0 9.432 0.024 9.648 ;
			RECT 0.0 9.672 0.024 9.888 ;
			RECT 0.0 9.912 0.024 10.128 ;
			RECT 0.0 10.152 0.024 10.368 ;
			RECT 0.0 10.392 0.024 10.608 ;
			RECT 0.0 10.632 0.024 10.848 ;
			RECT 0.0 10.872 0.024 11.088 ;
			RECT 0.0 11.112 0.024 11.328 ;
			RECT 0.0 11.352 0.024 11.568 ;
			RECT 0.0 11.592 0.024 11.808 ;
			RECT 0.0 11.832 0.024 12.048 ;
			RECT 0.0 12.072 0.024 12.288 ;
			RECT 0.0 12.312 0.024 12.528 ;
			RECT 0.0 12.552 0.024 12.768 ;
			RECT 0.0 12.792 0.024 13.008 ;
			RECT 0.0 13.032 0.024 13.248 ;
			RECT 0.0 13.272 0.024 13.488 ;
			RECT 0.0 13.512 0.024 13.728 ;
			RECT 0.0 13.752 0.024 13.968 ;
			RECT 0.0 13.992 0.024 14.208 ;
			RECT 0.0 14.232 0.024 14.448 ;
			RECT 0.0 14.472 0.024 14.688 ;
			RECT 0.0 14.712 0.024 14.928 ;
			RECT 0.0 14.952 0.024 15.168 ;
			RECT 0.0 15.192 0.024 15.216 ;
			RECT 0.0 15.24 0.024 15.456 ;
			RECT 0.0 15.48 0.024 15.696 ;
			RECT 0.0 15.72 0.024 15.936 ;
			RECT 0.0 15.96 0.024 16.176 ;
			RECT 0.0 16.2 0.024 16.416 ;
			RECT 0.0 16.44 0.024 16.656 ;
			RECT 0.0 16.68 0.024 16.896 ;
			RECT 0.0 16.92 0.024 17.136 ;
			RECT 0.0 17.16 0.024 17.376 ;
			RECT 0.0 17.4 0.024 17.616 ;
			RECT 0.0 17.64 0.024 17.856 ;
			RECT 0.0 17.88 0.024 18.096 ;
			RECT 0.0 18.12 0.024 18.336 ;
			RECT 0.0 18.36 0.024 18.576 ;
			RECT 0.0 18.6 0.024 18.816 ;
			RECT 0.0 18.84 0.024 19.056 ;
			RECT 0.0 19.08 0.024 19.296 ;
			RECT 0.0 19.32 0.024 19.536 ;
			RECT 0.0 19.56 0.024 19.776 ;
			RECT 0.0 19.8 0.024 20.016 ;
			RECT 0.0 20.04 0.024 20.256 ;
			RECT 0.0 20.28 0.024 20.496 ;
			RECT 0.0 20.52 0.024 20.736 ;
			RECT 0.0 20.76 0.024 20.976 ;
			RECT 0.0 21.0 0.024 21.216 ;
			RECT 0.0 21.24 0.024 21.456 ;
			RECT 0.0 21.48 0.024 21.696 ;
			RECT 0.0 21.72 0.024 21.936 ;
			RECT 0.0 21.96 0.024 22.176 ;
			RECT 0.0 22.2 0.024 22.416 ;
			RECT 0.0 22.44 0.024 22.656 ;
			RECT 0.0 22.68 0.024 22.896 ;
			RECT 0.0 22.92 0.024 23.136 ;
			RECT 0.0 23.16 0.024 23.376 ;
			RECT 0.0 23.4 0.024 23.616 ;
			RECT 0.0 23.64 0.024 23.856 ;
			RECT 0.0 23.88 0.024 24.096 ;
			RECT 0.0 24.12 0.024 24.336 ;
			RECT 0.0 24.36 0.024 24.576 ;
			RECT 0.0 24.6 0.024 24.816 ;
			RECT 0.0 24.84 0.024 25.056 ;
			RECT 0.0 25.08 0.024 25.296 ;
			RECT 0.0 25.32 0.024 25.536 ;
			RECT 0.0 25.56 0.024 25.776 ;
			RECT 0.0 25.8 0.024 26.016 ;
			RECT 0.0 26.04 0.024 26.256 ;
			RECT 0.0 26.28 0.024 26.496 ;
			RECT 0.0 26.52 0.024 26.736 ;
			RECT 0.0 26.76 0.024 26.976 ;
			RECT 0.0 27.0 0.024 27.216 ;
			RECT 0.0 27.24 0.024 27.456 ;
			RECT 0.0 27.48 0.024 27.696 ;
			RECT 0.0 27.72 0.024 27.936 ;
			RECT 0.0 27.96 0.024 28.176 ;
			RECT 0.0 28.2 0.024 28.416 ;
			RECT 0.0 28.44 0.024 28.656 ;
			RECT 0.0 28.68 0.024 28.896 ;
			RECT 0.0 28.92 0.024 29.136 ;
			RECT 0.0 29.16 0.024 29.376 ;
			RECT 0.0 29.4 0.024 29.616 ;
			RECT 0.0 29.64 0.024 29.856 ;
			RECT 0.0 29.88 0.024 30.096 ;
			RECT 0.0 30.12 0.024 30.336 ;
			RECT 0.0 30.36 0.024 30.384 ;
			RECT 0.0 30.408 0.024 30.624 ;
			RECT 0.0 30.648 0.024 30.864 ;
			RECT 0.0 30.888 0.024 31.104 ;
			RECT 0.0 31.128 0.024 31.344 ;
			RECT 0.0 31.368 0.024 31.584 ;
			RECT 0.0 31.608 0.024 31.824 ;
			RECT 0.0 31.848 0.024 32.064 ;
			RECT 0.0 32.088 0.024 32.304 ;
			RECT 0.0 32.328 0.024 32.544 ;
			RECT 0.0 32.568 0.024 32.784 ;
			RECT 0.0 32.808 0.024 33.024 ;
			RECT 0.0 33.048 0.024 33.264 ;
			RECT 0.0 33.288 0.024 33.504 ;
			RECT 0.0 33.528 0.024 33.744 ;
			RECT 0.0 33.768 0.024 33.984 ;
			RECT 0.0 34.008 0.024 34.224 ;
			RECT 0.0 34.248 0.024 34.464 ;
			RECT 0.0 34.488 0.024 34.704 ;
			RECT 0.0 34.728 0.024 34.944 ;
			RECT 0.0 34.968 0.024 35.184 ;
			RECT 0.0 35.208 0.024 35.424 ;
			RECT 0.0 35.448 0.024 35.664 ;
			RECT 0.0 35.688 0.024 35.904 ;
			RECT 0.0 35.928 0.024 36.144 ;
			RECT 0.0 36.168 0.024 36.384 ;
			RECT 0.0 36.408 0.024 36.624 ;
			RECT 0.0 36.648 0.024 36.864 ;
			RECT 0.0 36.888 0.024 37.104 ;
			RECT 0.0 37.128 0.024 37.344 ;
			RECT 0.0 37.368 0.024 37.584 ;
			RECT 0.0 37.608 0.024 37.824 ;
			RECT 0.0 37.848 0.024 38.064 ;
			RECT 0.0 38.088 0.024 38.304 ;
			RECT 0.0 38.328 0.024 38.544 ;
			RECT 0.0 38.568 0.024 38.784 ;
			RECT 0.0 38.808 0.024 39.024 ;
			RECT 0.0 39.048 0.024 39.264 ;
			RECT 0.0 39.288 0.024 39.504 ;
			RECT 0.0 39.528 0.024 39.744 ;
			RECT 0.0 39.768 0.024 39.984 ;
			RECT 0.0 40.008 0.024 40.224 ;
			RECT 0.0 40.248 0.024 40.464 ;
			RECT 0.0 40.488 0.024 40.704 ;
			RECT 0.0 40.728 0.024 40.944 ;
			RECT 0.0 40.968 0.024 41.184 ;
			RECT 0.0 41.208 0.024 41.424 ;
			RECT 0.0 41.448 0.024 41.664 ;
			RECT 0.0 41.688 0.024 41.904 ;
			RECT 0.0 41.928 0.024 42.144 ;
			RECT 0.0 42.168 0.024 42.384 ;
			RECT 0.0 42.408 0.024 42.624 ;
			RECT 0.0 42.648 0.024 42.864 ;
			RECT 0.0 42.888 0.024 43.104 ;
			RECT 0.0 43.128 0.024 43.344 ;
			RECT 0.0 43.368 0.024 43.584 ;
			RECT 0.0 43.608 0.024 43.824 ;
			RECT 0.0 43.848 0.024 44.064 ;
			RECT 0.0 44.088 0.024 44.304 ;
			RECT 0.0 44.328 0.024 44.544 ;
			RECT 0.0 44.568 0.024 44.784 ;
			RECT 0.0 44.808 0.024 45.024 ;
			RECT 0.0 45.048 0.024 45.264 ;
			RECT 0.0 45.288 0.024 45.504 ;
			RECT 0.0 45.528 0.024 45.552 ;
			RECT 0.0 45.576 0.024 45.792 ;
			RECT 0.0 45.816 0.024 46.032 ;
			RECT 0.0 46.056 0.024 46.272 ;
			RECT 0.0 46.296 0.024 46.512 ;
			RECT 0.0 46.536 0.024 46.752 ;
			RECT 0.0 46.776 0.024 46.992 ;
			RECT 0.0 47.016 0.024 47.232 ;
			RECT 0.0 47.256 0.024 47.28 ;
			RECT 0.0 47.304 0.024 47.52 ;
			RECT 0.0 47.544 0.024 47.76 ;
			RECT 0.0 33.6 0.024 47.784 ;

	END

END sram_asap7_64x256_1rw

MACRO sram_asap7_64x64_1rw
	CLASS BLOCK ;
	FOREIGN sram_asap7_64x64_1rw 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 8.36 BY 16.8 ;
	SYMMETRY X Y ;
	PIN clk
		DIRECTION INPUT ;
		USE CLOCK ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.408 0.024 15.432 ;

		END 

	END clk
	PIN rd_out[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.096 0.024 6.12 ;

		END 

	END rd_out[63]
	PIN rd_out[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.0 0.024 6.024 ;

		END 

	END rd_out[62]
	PIN rd_out[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.904 0.024 5.928 ;

		END 

	END rd_out[61]
	PIN rd_out[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.808 0.024 5.832 ;

		END 

	END rd_out[60]
	PIN rd_out[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.712 0.024 5.736 ;

		END 

	END rd_out[59]
	PIN rd_out[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.616 0.024 5.64 ;

		END 

	END rd_out[58]
	PIN rd_out[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.52 0.024 5.544 ;

		END 

	END rd_out[57]
	PIN rd_out[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.424 0.024 5.448 ;

		END 

	END rd_out[56]
	PIN rd_out[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.328 0.024 5.352 ;

		END 

	END rd_out[55]
	PIN rd_out[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.232 0.024 5.256 ;

		END 

	END rd_out[54]
	PIN rd_out[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.136 0.024 5.16 ;

		END 

	END rd_out[53]
	PIN rd_out[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 5.04 0.024 5.064 ;

		END 

	END rd_out[52]
	PIN rd_out[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.944 0.024 4.968 ;

		END 

	END rd_out[51]
	PIN rd_out[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.848 0.024 4.872 ;

		END 

	END rd_out[50]
	PIN rd_out[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.752 0.024 4.776 ;

		END 

	END rd_out[49]
	PIN rd_out[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.656 0.024 4.68 ;

		END 

	END rd_out[48]
	PIN rd_out[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.56 0.024 4.584 ;

		END 

	END rd_out[47]
	PIN rd_out[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.464 0.024 4.488 ;

		END 

	END rd_out[46]
	PIN rd_out[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.368 0.024 4.392 ;

		END 

	END rd_out[45]
	PIN rd_out[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.272 0.024 4.296 ;

		END 

	END rd_out[44]
	PIN rd_out[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.176 0.024 4.2 ;

		END 

	END rd_out[43]
	PIN rd_out[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 4.08 0.024 4.104 ;

		END 

	END rd_out[42]
	PIN rd_out[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.984 0.024 4.008 ;

		END 

	END rd_out[41]
	PIN rd_out[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.888 0.024 3.912 ;

		END 

	END rd_out[40]
	PIN rd_out[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.792 0.024 3.816 ;

		END 

	END rd_out[39]
	PIN rd_out[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.696 0.024 3.72 ;

		END 

	END rd_out[38]
	PIN rd_out[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.6 0.024 3.624 ;

		END 

	END rd_out[37]
	PIN rd_out[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.504 0.024 3.528 ;

		END 

	END rd_out[36]
	PIN rd_out[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.408 0.024 3.432 ;

		END 

	END rd_out[35]
	PIN rd_out[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.312 0.024 3.336 ;

		END 

	END rd_out[34]
	PIN rd_out[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.216 0.024 3.24 ;

		END 

	END rd_out[33]
	PIN rd_out[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.12 0.024 3.144 ;

		END 

	END rd_out[32]
	PIN rd_out[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 3.024 0.024 3.048 ;

		END 

	END rd_out[31]
	PIN rd_out[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.928 0.024 2.952 ;

		END 

	END rd_out[30]
	PIN rd_out[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.832 0.024 2.856 ;

		END 

	END rd_out[29]
	PIN rd_out[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.736 0.024 2.76 ;

		END 

	END rd_out[28]
	PIN rd_out[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.64 0.024 2.664 ;

		END 

	END rd_out[27]
	PIN rd_out[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.544 0.024 2.568 ;

		END 

	END rd_out[26]
	PIN rd_out[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.448 0.024 2.472 ;

		END 

	END rd_out[25]
	PIN rd_out[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.352 0.024 2.376 ;

		END 

	END rd_out[24]
	PIN rd_out[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.256 0.024 2.28 ;

		END 

	END rd_out[23]
	PIN rd_out[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.16 0.024 2.184 ;

		END 

	END rd_out[22]
	PIN rd_out[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 2.064 0.024 2.088 ;

		END 

	END rd_out[21]
	PIN rd_out[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.968 0.024 1.992 ;

		END 

	END rd_out[20]
	PIN rd_out[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.872 0.024 1.896 ;

		END 

	END rd_out[19]
	PIN rd_out[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.776 0.024 1.8 ;

		END 

	END rd_out[18]
	PIN rd_out[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.68 0.024 1.704 ;

		END 

	END rd_out[17]
	PIN rd_out[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.584 0.024 1.608 ;

		END 

	END rd_out[16]
	PIN rd_out[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.488 0.024 1.512 ;

		END 

	END rd_out[15]
	PIN rd_out[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.392 0.024 1.416 ;

		END 

	END rd_out[14]
	PIN rd_out[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.296 0.024 1.32 ;

		END 

	END rd_out[13]
	PIN rd_out[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.2 0.024 1.224 ;

		END 

	END rd_out[12]
	PIN rd_out[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.104 0.024 1.128 ;

		END 

	END rd_out[11]
	PIN rd_out[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 1.008 0.024 1.032 ;

		END 

	END rd_out[10]
	PIN rd_out[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.912 0.024 0.936 ;

		END 

	END rd_out[9]
	PIN rd_out[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.816 0.024 0.84 ;

		END 

	END rd_out[8]
	PIN rd_out[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.72 0.024 0.744 ;

		END 

	END rd_out[7]
	PIN rd_out[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.624 0.024 0.648 ;

		END 

	END rd_out[6]
	PIN rd_out[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.528 0.024 0.552 ;

		END 

	END rd_out[5]
	PIN rd_out[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.432 0.024 0.456 ;

		END 

	END rd_out[4]
	PIN rd_out[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.336 0.024 0.36 ;

		END 

	END rd_out[3]
	PIN rd_out[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.24 0.024 0.264 ;

		END 

	END rd_out[2]
	PIN rd_out[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.144 0.024 0.168 ;

		END 

	END rd_out[1]
	PIN rd_out[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 0.048 0.024 0.072 ;

		END 

	END rd_out[0]
	PIN we_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.216 0.024 15.24 ;

		END 

	END we_in
	PIN ce_in
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 15.312 0.024 15.336 ;

		END 

	END ce_in
	PIN addr_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.352 0.024 14.376 ;

		END 

	END addr_in[5]
	PIN addr_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.256 0.024 14.28 ;

		END 

	END addr_in[4]
	PIN addr_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.16 0.024 14.184 ;

		END 

	END addr_in[3]
	PIN addr_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 14.064 0.024 14.088 ;

		END 

	END addr_in[2]
	PIN addr_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.968 0.024 13.992 ;

		END 

	END addr_in[1]
	PIN addr_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.872 0.024 13.896 ;

		END 

	END addr_in[0]
	PIN wd_in[63]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 13.008 0.024 13.032 ;

		END 

	END wd_in[63]
	PIN wd_in[62]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.912 0.024 12.936 ;

		END 

	END wd_in[62]
	PIN wd_in[61]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.816 0.024 12.84 ;

		END 

	END wd_in[61]
	PIN wd_in[60]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.72 0.024 12.744 ;

		END 

	END wd_in[60]
	PIN wd_in[59]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.624 0.024 12.648 ;

		END 

	END wd_in[59]
	PIN wd_in[58]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.528 0.024 12.552 ;

		END 

	END wd_in[58]
	PIN wd_in[57]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.432 0.024 12.456 ;

		END 

	END wd_in[57]
	PIN wd_in[56]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.336 0.024 12.36 ;

		END 

	END wd_in[56]
	PIN wd_in[55]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.24 0.024 12.264 ;

		END 

	END wd_in[55]
	PIN wd_in[54]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.144 0.024 12.168 ;

		END 

	END wd_in[54]
	PIN wd_in[53]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 12.048 0.024 12.072 ;

		END 

	END wd_in[53]
	PIN wd_in[52]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.952 0.024 11.976 ;

		END 

	END wd_in[52]
	PIN wd_in[51]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.856 0.024 11.88 ;

		END 

	END wd_in[51]
	PIN wd_in[50]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.76 0.024 11.784 ;

		END 

	END wd_in[50]
	PIN wd_in[49]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.664 0.024 11.688 ;

		END 

	END wd_in[49]
	PIN wd_in[48]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.568 0.024 11.592 ;

		END 

	END wd_in[48]
	PIN wd_in[47]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.472 0.024 11.496 ;

		END 

	END wd_in[47]
	PIN wd_in[46]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.376 0.024 11.4 ;

		END 

	END wd_in[46]
	PIN wd_in[45]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.28 0.024 11.304 ;

		END 

	END wd_in[45]
	PIN wd_in[44]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.184 0.024 11.208 ;

		END 

	END wd_in[44]
	PIN wd_in[43]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 11.088 0.024 11.112 ;

		END 

	END wd_in[43]
	PIN wd_in[42]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.992 0.024 11.016 ;

		END 

	END wd_in[42]
	PIN wd_in[41]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.896 0.024 10.92 ;

		END 

	END wd_in[41]
	PIN wd_in[40]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.8 0.024 10.824 ;

		END 

	END wd_in[40]
	PIN wd_in[39]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.704 0.024 10.728 ;

		END 

	END wd_in[39]
	PIN wd_in[38]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.608 0.024 10.632 ;

		END 

	END wd_in[38]
	PIN wd_in[37]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.512 0.024 10.536 ;

		END 

	END wd_in[37]
	PIN wd_in[36]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.416 0.024 10.44 ;

		END 

	END wd_in[36]
	PIN wd_in[35]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.32 0.024 10.344 ;

		END 

	END wd_in[35]
	PIN wd_in[34]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.224 0.024 10.248 ;

		END 

	END wd_in[34]
	PIN wd_in[33]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.128 0.024 10.152 ;

		END 

	END wd_in[33]
	PIN wd_in[32]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 10.032 0.024 10.056 ;

		END 

	END wd_in[32]
	PIN wd_in[31]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.936 0.024 9.96 ;

		END 

	END wd_in[31]
	PIN wd_in[30]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.84 0.024 9.864 ;

		END 

	END wd_in[30]
	PIN wd_in[29]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.744 0.024 9.768 ;

		END 

	END wd_in[29]
	PIN wd_in[28]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.648 0.024 9.672 ;

		END 

	END wd_in[28]
	PIN wd_in[27]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.552 0.024 9.576 ;

		END 

	END wd_in[27]
	PIN wd_in[26]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.456 0.024 9.48 ;

		END 

	END wd_in[26]
	PIN wd_in[25]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.36 0.024 9.384 ;

		END 

	END wd_in[25]
	PIN wd_in[24]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.264 0.024 9.288 ;

		END 

	END wd_in[24]
	PIN wd_in[23]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.168 0.024 9.192 ;

		END 

	END wd_in[23]
	PIN wd_in[22]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 9.072 0.024 9.096 ;

		END 

	END wd_in[22]
	PIN wd_in[21]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.976 0.024 9.0 ;

		END 

	END wd_in[21]
	PIN wd_in[20]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.88 0.024 8.904 ;

		END 

	END wd_in[20]
	PIN wd_in[19]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.784 0.024 8.808 ;

		END 

	END wd_in[19]
	PIN wd_in[18]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.688 0.024 8.712 ;

		END 

	END wd_in[18]
	PIN wd_in[17]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.592 0.024 8.616 ;

		END 

	END wd_in[17]
	PIN wd_in[16]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.496 0.024 8.52 ;

		END 

	END wd_in[16]
	PIN wd_in[15]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.4 0.024 8.424 ;

		END 

	END wd_in[15]
	PIN wd_in[14]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.304 0.024 8.328 ;

		END 

	END wd_in[14]
	PIN wd_in[13]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.208 0.024 8.232 ;

		END 

	END wd_in[13]
	PIN wd_in[12]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.112 0.024 8.136 ;

		END 

	END wd_in[12]
	PIN wd_in[11]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 8.016 0.024 8.04 ;

		END 

	END wd_in[11]
	PIN wd_in[10]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.92 0.024 7.944 ;

		END 

	END wd_in[10]
	PIN wd_in[9]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.824 0.024 7.848 ;

		END 

	END wd_in[9]
	PIN wd_in[8]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.728 0.024 7.752 ;

		END 

	END wd_in[8]
	PIN wd_in[7]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.632 0.024 7.656 ;

		END 

	END wd_in[7]
	PIN wd_in[6]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.536 0.024 7.56 ;

		END 

	END wd_in[6]
	PIN wd_in[5]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.44 0.024 7.464 ;

		END 

	END wd_in[5]
	PIN wd_in[4]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.344 0.024 7.368 ;

		END 

	END wd_in[4]
	PIN wd_in[3]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.248 0.024 7.272 ;

		END 

	END wd_in[3]
	PIN wd_in[2]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.152 0.024 7.176 ;

		END 

	END wd_in[2]
	PIN wd_in[1]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 7.056 0.024 7.08 ;

		END 

	END wd_in[1]
	PIN wd_in[0]
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER M4 ;
			RECT 0.0 6.96 0.024 6.984 ;

		END 

	END wd_in[0]
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.0 8.312 0.096 ;
			RECT 0.048 0.768 8.312 0.864 ;
			RECT 0.048 1.536 8.312 1.632 ;
			RECT 0.048 2.304 8.312 2.4 ;
			RECT 0.048 3.072 8.312 3.168 ;
			RECT 0.048 3.84 8.312 3.936 ;
			RECT 0.048 4.608 8.312 4.704 ;
			RECT 0.048 5.376 8.312 5.472 ;
			RECT 0.048 6.144 8.312 6.24 ;
			RECT 0.048 6.912 8.312 7.008 ;
			RECT 0.048 7.68 8.312 7.776 ;
			RECT 0.048 8.448 8.312 8.544 ;
			RECT 0.048 9.216 8.312 9.312 ;
			RECT 0.048 9.984 8.312 10.08 ;
			RECT 0.048 10.752 8.312 10.848 ;
			RECT 0.048 11.52 8.312 11.616 ;
			RECT 0.048 12.288 8.312 12.384 ;
			RECT 0.048 13.056 8.312 13.152 ;
			RECT 0.048 13.824 8.312 13.92 ;
			RECT 0.048 14.592 8.312 14.688 ;
			RECT 0.048 15.36 8.312 15.456 ;
			RECT 0.048 16.128 8.312 16.224 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT 
			LAYER M4 ;
			RECT 0.048 0.384 8.312 0.48 ;
			RECT 0.048 1.152 8.312 1.248 ;
			RECT 0.048 1.92 8.312 2.016 ;
			RECT 0.048 2.688 8.312 2.784 ;
			RECT 0.048 3.456 8.312 3.552 ;
			RECT 0.048 4.224 8.312 4.32 ;
			RECT 0.048 4.992 8.312 5.088 ;
			RECT 0.048 5.76 8.312 5.856 ;
			RECT 0.048 6.528 8.312 6.624 ;
			RECT 0.048 7.296 8.312 7.392 ;
			RECT 0.048 8.064 8.312 8.16 ;
			RECT 0.048 8.832 8.312 8.928 ;
			RECT 0.048 9.6 8.312 9.696 ;
			RECT 0.048 10.368 8.312 10.464 ;
			RECT 0.048 11.136 8.312 11.232 ;
			RECT 0.048 11.904 8.312 12.0 ;
			RECT 0.048 12.672 8.312 12.768 ;
			RECT 0.048 13.44 8.312 13.536 ;
			RECT 0.048 14.208 8.312 14.304 ;
			RECT 0.048 14.976 8.312 15.072 ;
			RECT 0.048 15.744 8.312 15.84 ;
			RECT 0.048 16.512 8.312 16.608 ;

		END 

	END VDD
	OBS
			LAYER M1 ;
			RECT 0.0 0.0 8.36 16.8 ;
			LAYER M2 ;
			RECT 0.0 0.0 8.36 16.8 ;
			LAYER M3 ;
			RECT 0.0 0.0 8.36 16.8 ;
			LAYER M4 ;
			RECT 0.024 0.0 0.048 16.8 ;
			RECT 8.312 0.0 8.36 16.8 ;
			RECT 0.048 0.0 8.312 0.0 ;
			RECT 0.048 0.096 8.312 0.384 ;
			RECT 0.048 0.48 8.312 0.768 ;
			RECT 0.048 0.864 8.312 1.152 ;
			RECT 0.048 1.248 8.312 1.536 ;
			RECT 0.048 1.632 8.312 1.92 ;
			RECT 0.048 2.016 8.312 2.304 ;
			RECT 0.048 2.4 8.312 2.688 ;
			RECT 0.048 2.784 8.312 3.072 ;
			RECT 0.048 3.168 8.312 3.456 ;
			RECT 0.048 3.552 8.312 3.84 ;
			RECT 0.048 3.936 8.312 4.224 ;
			RECT 0.048 4.32 8.312 4.608 ;
			RECT 0.048 4.704 8.312 4.992 ;
			RECT 0.048 5.088 8.312 5.376 ;
			RECT 0.048 5.472 8.312 5.76 ;
			RECT 0.048 5.856 8.312 6.144 ;
			RECT 0.048 6.24 8.312 6.528 ;
			RECT 0.048 6.624 8.312 6.912 ;
			RECT 0.048 7.008 8.312 7.296 ;
			RECT 0.048 7.392 8.312 7.68 ;
			RECT 0.048 7.776 8.312 8.064 ;
			RECT 0.048 8.16 8.312 8.448 ;
			RECT 0.048 8.544 8.312 8.832 ;
			RECT 0.048 8.928 8.312 9.216 ;
			RECT 0.048 9.312 8.312 9.6 ;
			RECT 0.048 9.696 8.312 9.984 ;
			RECT 0.048 10.08 8.312 10.368 ;
			RECT 0.048 10.464 8.312 10.752 ;
			RECT 0.048 10.848 8.312 11.136 ;
			RECT 0.048 11.232 8.312 11.52 ;
			RECT 0.048 11.616 8.312 11.904 ;
			RECT 0.048 12.0 8.312 12.288 ;
			RECT 0.048 12.384 8.312 12.672 ;
			RECT 0.048 12.768 8.312 13.056 ;
			RECT 0.048 13.152 8.312 13.44 ;
			RECT 0.048 13.536 8.312 13.824 ;
			RECT 0.048 13.92 8.312 14.208 ;
			RECT 0.048 14.304 8.312 14.592 ;
			RECT 0.048 14.688 8.312 14.976 ;
			RECT 0.048 15.072 8.312 15.36 ;
			RECT 0.048 15.456 8.312 15.744 ;
			RECT 0.048 15.84 8.312 16.128 ;
			RECT 0.048 16.224 8.312 16.512 ;
			RECT 0.048 16.608 8.312 16.8 ;
			RECT 0.0 0.0 0.024 0.048 ;
			RECT 0.0 0.072 0.024 0.144 ;
			RECT 0.0 0.168 0.024 0.24 ;
			RECT 0.0 0.264 0.024 0.336 ;
			RECT 0.0 0.36 0.024 0.432 ;
			RECT 0.0 0.456 0.024 0.528 ;
			RECT 0.0 0.552 0.024 0.624 ;
			RECT 0.0 0.648 0.024 0.72 ;
			RECT 0.0 0.744 0.024 0.816 ;
			RECT 0.0 0.84 0.024 0.912 ;
			RECT 0.0 0.936 0.024 1.008 ;
			RECT 0.0 1.032 0.024 1.104 ;
			RECT 0.0 1.128 0.024 1.2 ;
			RECT 0.0 1.224 0.024 1.296 ;
			RECT 0.0 1.32 0.024 1.392 ;
			RECT 0.0 1.416 0.024 1.488 ;
			RECT 0.0 1.512 0.024 1.584 ;
			RECT 0.0 1.608 0.024 1.68 ;
			RECT 0.0 1.704 0.024 1.776 ;
			RECT 0.0 1.8 0.024 1.872 ;
			RECT 0.0 1.896 0.024 1.968 ;
			RECT 0.0 1.992 0.024 2.064 ;
			RECT 0.0 2.088 0.024 2.16 ;
			RECT 0.0 2.184 0.024 2.256 ;
			RECT 0.0 2.28 0.024 2.352 ;
			RECT 0.0 2.376 0.024 2.448 ;
			RECT 0.0 2.472 0.024 2.544 ;
			RECT 0.0 2.568 0.024 2.64 ;
			RECT 0.0 2.664 0.024 2.736 ;
			RECT 0.0 2.76 0.024 2.832 ;
			RECT 0.0 2.856 0.024 2.928 ;
			RECT 0.0 2.952 0.024 3.024 ;
			RECT 0.0 3.048 0.024 3.12 ;
			RECT 0.0 3.144 0.024 3.216 ;
			RECT 0.0 3.24 0.024 3.312 ;
			RECT 0.0 3.336 0.024 3.408 ;
			RECT 0.0 3.432 0.024 3.504 ;
			RECT 0.0 3.528 0.024 3.6 ;
			RECT 0.0 3.624 0.024 3.696 ;
			RECT 0.0 3.72 0.024 3.792 ;
			RECT 0.0 3.816 0.024 3.888 ;
			RECT 0.0 3.912 0.024 3.984 ;
			RECT 0.0 4.008 0.024 4.08 ;
			RECT 0.0 4.104 0.024 4.176 ;
			RECT 0.0 4.2 0.024 4.272 ;
			RECT 0.0 4.296 0.024 4.368 ;
			RECT 0.0 4.392 0.024 4.464 ;
			RECT 0.0 4.488 0.024 4.56 ;
			RECT 0.0 4.584 0.024 4.656 ;
			RECT 0.0 4.68 0.024 4.752 ;
			RECT 0.0 4.776 0.024 4.848 ;
			RECT 0.0 4.872 0.024 4.944 ;
			RECT 0.0 4.968 0.024 5.04 ;
			RECT 0.0 5.064 0.024 5.136 ;
			RECT 0.0 5.16 0.024 5.232 ;
			RECT 0.0 5.256 0.024 5.328 ;
			RECT 0.0 5.352 0.024 5.424 ;
			RECT 0.0 5.448 0.024 5.52 ;
			RECT 0.0 5.544 0.024 5.616 ;
			RECT 0.0 5.64 0.024 5.712 ;
			RECT 0.0 5.736 0.024 5.808 ;
			RECT 0.0 5.832 0.024 5.904 ;
			RECT 0.0 5.928 0.024 6.0 ;
			RECT 0.0 6.024 0.024 6.096 ;
			RECT 0.0 6.12 0.024 6.96 ;
			RECT 0.0 6.984 0.024 7.056 ;
			RECT 0.0 7.08 0.024 7.152 ;
			RECT 0.0 7.176 0.024 7.248 ;
			RECT 0.0 7.272 0.024 7.344 ;
			RECT 0.0 7.368 0.024 7.44 ;
			RECT 0.0 7.464 0.024 7.536 ;
			RECT 0.0 7.56 0.024 7.632 ;
			RECT 0.0 7.656 0.024 7.728 ;
			RECT 0.0 7.752 0.024 7.824 ;
			RECT 0.0 7.848 0.024 7.92 ;
			RECT 0.0 7.944 0.024 8.016 ;
			RECT 0.0 8.04 0.024 8.112 ;
			RECT 0.0 8.136 0.024 8.208 ;
			RECT 0.0 8.232 0.024 8.304 ;
			RECT 0.0 8.328 0.024 8.4 ;
			RECT 0.0 8.424 0.024 8.496 ;
			RECT 0.0 8.52 0.024 8.592 ;
			RECT 0.0 8.616 0.024 8.688 ;
			RECT 0.0 8.712 0.024 8.784 ;
			RECT 0.0 8.808 0.024 8.88 ;
			RECT 0.0 8.904 0.024 8.976 ;
			RECT 0.0 9.0 0.024 9.072 ;
			RECT 0.0 9.096 0.024 9.168 ;
			RECT 0.0 9.192 0.024 9.264 ;
			RECT 0.0 9.288 0.024 9.36 ;
			RECT 0.0 9.384 0.024 9.456 ;
			RECT 0.0 9.48 0.024 9.552 ;
			RECT 0.0 9.576 0.024 9.648 ;
			RECT 0.0 9.672 0.024 9.744 ;
			RECT 0.0 9.768 0.024 9.84 ;
			RECT 0.0 9.864 0.024 9.936 ;
			RECT 0.0 9.96 0.024 10.032 ;
			RECT 0.0 10.056 0.024 10.128 ;
			RECT 0.0 10.152 0.024 10.224 ;
			RECT 0.0 10.248 0.024 10.32 ;
			RECT 0.0 10.344 0.024 10.416 ;
			RECT 0.0 10.44 0.024 10.512 ;
			RECT 0.0 10.536 0.024 10.608 ;
			RECT 0.0 10.632 0.024 10.704 ;
			RECT 0.0 10.728 0.024 10.8 ;
			RECT 0.0 10.824 0.024 10.896 ;
			RECT 0.0 10.92 0.024 10.992 ;
			RECT 0.0 11.016 0.024 11.088 ;
			RECT 0.0 11.112 0.024 11.184 ;
			RECT 0.0 11.208 0.024 11.28 ;
			RECT 0.0 11.304 0.024 11.376 ;
			RECT 0.0 11.4 0.024 11.472 ;
			RECT 0.0 11.496 0.024 11.568 ;
			RECT 0.0 11.592 0.024 11.664 ;
			RECT 0.0 11.688 0.024 11.76 ;
			RECT 0.0 11.784 0.024 11.856 ;
			RECT 0.0 11.88 0.024 11.952 ;
			RECT 0.0 11.976 0.024 12.048 ;
			RECT 0.0 12.072 0.024 12.144 ;
			RECT 0.0 12.168 0.024 12.24 ;
			RECT 0.0 12.264 0.024 12.336 ;
			RECT 0.0 12.36 0.024 12.432 ;
			RECT 0.0 12.456 0.024 12.528 ;
			RECT 0.0 12.552 0.024 12.624 ;
			RECT 0.0 12.648 0.024 12.72 ;
			RECT 0.0 12.744 0.024 12.816 ;
			RECT 0.0 12.84 0.024 12.912 ;
			RECT 0.0 12.936 0.024 13.008 ;
			RECT 0.0 13.032 0.024 13.872 ;
			RECT 0.0 13.896 0.024 13.968 ;
			RECT 0.0 13.992 0.024 14.064 ;
			RECT 0.0 14.088 0.024 14.16 ;
			RECT 0.0 14.184 0.024 14.256 ;
			RECT 0.0 14.28 0.024 14.352 ;
			RECT 0.0 14.376 0.024 14.448 ;
			RECT 0.0 14.472 0.024 14.544 ;
			RECT 0.0 14.568 0.024 14.64 ;
			RECT 0.0 14.664 0.024 14.736 ;
			RECT 0.0 14.76 0.024 14.832 ;
			RECT 0.0 14.856 0.024 14.928 ;
			RECT 0.0 14.952 0.024 15.024 ;
			RECT 0.0 15.048 0.024 15.12 ;
			RECT 0.0 15.144 0.024 15.216 ;
			RECT 0.0 15.24 0.024 15.312 ;
			RECT 0.0 15.336 0.024 15.408 ;
			RECT 0.0 15.432 0.024 15.504 ;
			RECT 0.0 15.528 0.024 15.6 ;
			RECT 0.0 15.624 0.024 15.696 ;
			RECT 0.0 15.72 0.024 15.792 ;
			RECT 0.0 15.816 0.024 15.888 ;
			RECT 0.0 15.912 0.024 15.984 ;
			RECT 0.0 16.008 0.024 16.08 ;
			RECT 0.0 16.104 0.024 16.176 ;
			RECT 0.0 16.2 0.024 16.272 ;
			RECT 0.0 16.296 0.024 16.368 ;
			RECT 0.0 16.392 0.024 16.464 ;
			RECT 0.0 16.488 0.024 16.56 ;
			RECT 0.0 16.584 0.024 16.656 ;
			RECT 0.0 16.68 0.024 16.752 ;
			RECT 0.0 16.776 0.024 16.848 ;
			RECT 0.0 16.872 0.024 16.944 ;
			RECT 0.0 16.968 0.024 17.04 ;
			RECT 0.0 17.064 0.024 17.136 ;
			RECT 0.0 17.16 0.024 17.232 ;
			RECT 0.0 17.256 0.024 17.328 ;
			RECT 0.0 17.352 0.024 17.424 ;
			RECT 0.0 17.448 0.024 17.52 ;
			RECT 0.0 17.544 0.024 17.616 ;
			RECT 0.0 17.64 0.024 17.712 ;
			RECT 0.0 17.736 0.024 17.808 ;
			RECT 0.0 17.832 0.024 17.904 ;
			RECT 0.0 17.928 0.024 18.0 ;
			RECT 0.0 18.024 0.024 18.096 ;
			RECT 0.0 18.12 0.024 18.192 ;
			RECT 0.0 18.216 0.024 18.288 ;
			RECT 0.0 18.312 0.024 18.384 ;
			RECT 0.0 18.408 0.024 18.48 ;
			RECT 0.0 18.504 0.024 18.576 ;
			RECT 0.0 18.6 0.024 18.672 ;
			RECT 0.0 18.696 0.024 18.768 ;
			RECT 0.0 18.792 0.024 18.864 ;
			RECT 0.0 18.888 0.024 18.96 ;
			RECT 0.0 18.984 0.024 19.056 ;
			RECT 0.0 19.08 0.024 19.152 ;
			RECT 0.0 19.176 0.024 19.248 ;
			RECT 0.0 19.272 0.024 19.344 ;
			RECT 0.0 19.368 0.024 19.44 ;
			RECT 0.0 19.464 0.024 19.536 ;
			RECT 0.0 19.56 0.024 19.632 ;
			RECT 0.0 19.656 0.024 19.728 ;
			RECT 0.0 19.752 0.024 19.824 ;
			RECT 0.0 19.848 0.024 19.92 ;
			RECT 0.0 19.944 0.024 20.784 ;
			RECT 0.0 20.808 0.024 20.88 ;
			RECT 0.0 20.904 0.024 20.976 ;
			RECT 0.0 21.0 0.024 21.072 ;
			RECT 0.0 21.096 0.024 21.168 ;
			RECT 0.0 21.192 0.024 21.264 ;
			RECT 0.0 21.288 0.024 22.128 ;
			RECT 0.0 22.152 0.024 22.224 ;
			RECT 0.0 22.248 0.024 22.32 ;
			RECT 0.0 16.8 0.024 22.344 ;

	END

END sram_asap7_64x64_1rw

END LIBRARY
